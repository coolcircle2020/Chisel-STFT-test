module ComplexAdd(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) + $signed(io_op2_re); // @[Butterfly.scala 21:13]
  assign io_res_im = $signed(io_op1_im) + $signed(io_op2_im); // @[Butterfly.scala 22:13]
endmodule
module ComplexSub(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  assign io_res_re = $signed(io_op1_re) - $signed(io_op2_re); // @[Butterfly.scala 35:13]
  assign io_res_im = $signed(io_op1_im) - $signed(io_op2_im); // @[Butterfly.scala 36:13]
endmodule
module ComplexMul(
  input  [31:0] io_op1_re,
  input  [31:0] io_op1_im,
  input  [31:0] io_op2_re,
  input  [31:0] io_op2_im,
  output [31:0] io_res_re,
  output [31:0] io_res_im
);
  wire [63:0] _T = $signed(io_op1_re) * $signed(io_op2_re); // @[Butterfly.scala 57:28]
  wire [63:0] _T_1 = $signed(io_op1_im) * $signed(io_op2_im); // @[Butterfly.scala 57:52]
  wire [63:0] _T_4 = $signed(_T) - $signed(_T_1); // @[Butterfly.scala 57:40]
  wire [63:0] _T_5 = $signed(io_op1_re) * $signed(io_op2_im); // @[Butterfly.scala 58:28]
  wire [63:0] _T_6 = $signed(io_op1_im) * $signed(io_op2_re); // @[Butterfly.scala 58:52]
  wire [63:0] _T_9 = $signed(_T_5) + $signed(_T_6); // @[Butterfly.scala 58:40]
  wire [47:0] _GEN_0 = _T_4[63:16]; // @[Butterfly.scala 57:15]
  wire [47:0] _GEN_2 = _T_9[63:16]; // @[Butterfly.scala 58:15]
  assign io_res_re = _GEN_0[31:0]; // @[Butterfly.scala 57:15]
  assign io_res_im = _GEN_2[31:0]; // @[Butterfly.scala 58:15]
endmodule
module Butterfly(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input  [31:0] io_wn_re,
  input  [31:0] io_wn_im,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexMul_io_op1_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op1_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_op2_im; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_re; // @[Butterfly.scala 63:22]
  wire [31:0] ComplexMul_io_res_im; // @[Butterfly.scala 63:22]
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  ComplexMul ComplexMul ( // @[Butterfly.scala 63:22]
    .io_op1_re(ComplexMul_io_op1_re),
    .io_op1_im(ComplexMul_io_op1_im),
    .io_op2_re(ComplexMul_io_op2_re),
    .io_op2_im(ComplexMul_io_op2_im),
    .io_res_re(ComplexMul_io_res_re),
    .io_res_im(ComplexMul_io_res_im)
  );
  assign io_out1_re = ComplexAdd_io_res_re; // @[Butterfly.scala 84:11]
  assign io_out1_im = ComplexAdd_io_res_im; // @[Butterfly.scala 84:11]
  assign io_out2_re = ComplexMul_io_res_re; // @[Butterfly.scala 85:11]
  assign io_out2_im = ComplexMul_io_res_im; // @[Butterfly.scala 85:11]
  assign ComplexAdd_io_op1_re = io_in1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = io_in1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = io_in2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = io_in2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = io_in1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = io_in1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = io_in2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = io_in2_im; // @[Butterfly.scala 42:17]
  assign ComplexMul_io_op1_re = ComplexSub_io_res_re; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op1_im = ComplexSub_io_res_im; // @[Butterfly.scala 64:17]
  assign ComplexMul_io_op2_re = io_wn_re; // @[Butterfly.scala 65:17]
  assign ComplexMul_io_op2_im = io_wn_im; // @[Butterfly.scala 65:17]
endmodule
module Switch(
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_sel,
  output [31:0] io_out1_re,
  output [31:0] io_out1_im,
  output [31:0] io_out2_re,
  output [31:0] io_out2_im
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[Butterfly.scala 105:11]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[Butterfly.scala 105:11]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[Butterfly.scala 106:11]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[Butterfly.scala 106:11]
endmodule
module FFT(
  input         clock,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut1_re,
  output [31:0] io_dOut1_im,
  output [31:0] io_dOut2_re,
  output [31:0] io_dOut2_im,
  output        io_dout_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [31:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [31:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [31:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [31:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [31:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [31:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [31:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [31:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [31:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [31:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [31:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [31:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [31:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [31:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [31:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [31:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [31:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [31:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [31:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [31:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [31:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [31:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [31:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [31:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [31:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [31:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [31:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [31:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [31:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [31:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [31:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [31:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [31:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [31:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [31:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [31:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [31:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [31:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [31:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [31:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [31:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [31:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [31:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [31:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [31:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [31:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [31:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [31:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [31:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [31:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [31:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [31:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [31:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [31:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [31:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [31:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [31:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [31:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [31:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [31:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [31:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [31:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [31:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [31:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [31:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [31:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [31:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [31:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [31:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [31:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [31:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [31:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [31:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [31:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [31:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [31:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [31:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [31:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [31:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [31:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [31:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [31:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [31:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [31:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [31:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [31:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [31:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [31:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [31:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [31:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [31:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [31:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [31:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [31:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [31:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [31:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [31:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [31:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [31:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [31:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [31:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [31:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [31:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [31:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [31:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [31:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [31:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [31:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [31:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [31:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [31:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [31:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [31:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [31:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [31:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [31:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [31:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [31:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [31:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [31:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [31:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [31:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [31:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [31:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [31:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [31:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [31:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [31:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [31:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [31:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [31:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [31:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [31:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [31:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [31:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [31:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [31:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [31:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [31:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [31:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [31:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [31:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [31:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [31:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [31:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [31:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [31:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [31:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [31:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [31:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [31:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [31:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [31:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [31:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [31:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [31:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [31:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [31:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [31:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [31:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [31:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [31:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [31:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [31:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [31:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [31:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [31:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [31:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [31:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [31:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [31:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [31:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [31:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [31:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [31:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [31:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [31:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [31:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [31:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [31:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [31:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [31:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [31:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [31:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [31:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [31:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [31:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [31:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [31:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [31:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [31:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [31:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [31:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [31:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [31:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [31:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [31:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [31:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [31:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [31:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [31:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [31:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [31:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [31:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [31:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [31:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [31:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [31:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [31:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [31:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [31:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [31:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [31:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [31:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [31:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [31:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [31:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [31:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [31:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [31:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [31:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [31:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [31:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [31:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [31:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [31:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [31:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [31:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [31:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [31:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [31:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [31:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [31:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [31:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [31:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [31:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [31:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [31:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [31:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [31:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [31:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [31:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [31:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [31:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [31:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [31:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [31:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [31:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [31:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [31:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [31:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [31:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
  reg [31:0] _RAND_2049;
  reg [31:0] _RAND_2050;
  reg [31:0] _RAND_2051;
  reg [31:0] _RAND_2052;
  reg [31:0] _RAND_2053;
  reg [31:0] _RAND_2054;
  reg [31:0] _RAND_2055;
  reg [31:0] _RAND_2056;
  reg [31:0] _RAND_2057;
  reg [31:0] _RAND_2058;
  reg [31:0] _RAND_2059;
  reg [31:0] _RAND_2060;
  reg [31:0] _RAND_2061;
  reg [31:0] _RAND_2062;
  reg [31:0] _RAND_2063;
  reg [31:0] _RAND_2064;
  reg [31:0] _RAND_2065;
  reg [31:0] _RAND_2066;
  reg [31:0] _RAND_2067;
  reg [31:0] _RAND_2068;
  reg [31:0] _RAND_2069;
  reg [31:0] _RAND_2070;
  reg [31:0] _RAND_2071;
  reg [31:0] _RAND_2072;
  reg [31:0] _RAND_2073;
  reg [31:0] _RAND_2074;
  reg [31:0] _RAND_2075;
  reg [31:0] _RAND_2076;
  reg [31:0] _RAND_2077;
  reg [31:0] _RAND_2078;
  reg [31:0] _RAND_2079;
  reg [31:0] _RAND_2080;
  reg [31:0] _RAND_2081;
  reg [31:0] _RAND_2082;
  reg [31:0] _RAND_2083;
  reg [31:0] _RAND_2084;
  reg [31:0] _RAND_2085;
  reg [31:0] _RAND_2086;
  reg [31:0] _RAND_2087;
  reg [31:0] _RAND_2088;
  reg [31:0] _RAND_2089;
  reg [31:0] _RAND_2090;
  reg [31:0] _RAND_2091;
  reg [31:0] _RAND_2092;
  reg [31:0] _RAND_2093;
  reg [31:0] _RAND_2094;
  reg [31:0] _RAND_2095;
  reg [31:0] _RAND_2096;
  reg [31:0] _RAND_2097;
  reg [31:0] _RAND_2098;
  reg [31:0] _RAND_2099;
  reg [31:0] _RAND_2100;
  reg [31:0] _RAND_2101;
  reg [31:0] _RAND_2102;
  reg [31:0] _RAND_2103;
  reg [31:0] _RAND_2104;
  reg [31:0] _RAND_2105;
  reg [31:0] _RAND_2106;
  reg [31:0] _RAND_2107;
  reg [31:0] _RAND_2108;
  reg [31:0] _RAND_2109;
  reg [31:0] _RAND_2110;
  reg [31:0] _RAND_2111;
  reg [31:0] _RAND_2112;
  reg [31:0] _RAND_2113;
  reg [31:0] _RAND_2114;
  reg [31:0] _RAND_2115;
  reg [31:0] _RAND_2116;
  reg [31:0] _RAND_2117;
  reg [31:0] _RAND_2118;
  reg [31:0] _RAND_2119;
  reg [31:0] _RAND_2120;
  reg [31:0] _RAND_2121;
  reg [31:0] _RAND_2122;
  reg [31:0] _RAND_2123;
  reg [31:0] _RAND_2124;
  reg [31:0] _RAND_2125;
  reg [31:0] _RAND_2126;
  reg [31:0] _RAND_2127;
  reg [31:0] _RAND_2128;
  reg [31:0] _RAND_2129;
  reg [31:0] _RAND_2130;
  reg [31:0] _RAND_2131;
  reg [31:0] _RAND_2132;
  reg [31:0] _RAND_2133;
  reg [31:0] _RAND_2134;
  reg [31:0] _RAND_2135;
  reg [31:0] _RAND_2136;
  reg [31:0] _RAND_2137;
  reg [31:0] _RAND_2138;
  reg [31:0] _RAND_2139;
  reg [31:0] _RAND_2140;
  reg [31:0] _RAND_2141;
  reg [31:0] _RAND_2142;
  reg [31:0] _RAND_2143;
  reg [31:0] _RAND_2144;
  reg [31:0] _RAND_2145;
  reg [31:0] _RAND_2146;
  reg [31:0] _RAND_2147;
  reg [31:0] _RAND_2148;
  reg [31:0] _RAND_2149;
  reg [31:0] _RAND_2150;
  reg [31:0] _RAND_2151;
  reg [31:0] _RAND_2152;
  reg [31:0] _RAND_2153;
  reg [31:0] _RAND_2154;
  reg [31:0] _RAND_2155;
  reg [31:0] _RAND_2156;
  reg [31:0] _RAND_2157;
  reg [31:0] _RAND_2158;
  reg [31:0] _RAND_2159;
  reg [31:0] _RAND_2160;
  reg [31:0] _RAND_2161;
  reg [31:0] _RAND_2162;
  reg [31:0] _RAND_2163;
  reg [31:0] _RAND_2164;
  reg [31:0] _RAND_2165;
  reg [31:0] _RAND_2166;
  reg [31:0] _RAND_2167;
  reg [31:0] _RAND_2168;
  reg [31:0] _RAND_2169;
  reg [31:0] _RAND_2170;
  reg [31:0] _RAND_2171;
  reg [31:0] _RAND_2172;
  reg [31:0] _RAND_2173;
  reg [31:0] _RAND_2174;
  reg [31:0] _RAND_2175;
  reg [31:0] _RAND_2176;
  reg [31:0] _RAND_2177;
  reg [31:0] _RAND_2178;
  reg [31:0] _RAND_2179;
  reg [31:0] _RAND_2180;
  reg [31:0] _RAND_2181;
  reg [31:0] _RAND_2182;
  reg [31:0] _RAND_2183;
  reg [31:0] _RAND_2184;
  reg [31:0] _RAND_2185;
  reg [31:0] _RAND_2186;
  reg [31:0] _RAND_2187;
  reg [31:0] _RAND_2188;
  reg [31:0] _RAND_2189;
  reg [31:0] _RAND_2190;
  reg [31:0] _RAND_2191;
  reg [31:0] _RAND_2192;
  reg [31:0] _RAND_2193;
  reg [31:0] _RAND_2194;
  reg [31:0] _RAND_2195;
  reg [31:0] _RAND_2196;
  reg [31:0] _RAND_2197;
  reg [31:0] _RAND_2198;
  reg [31:0] _RAND_2199;
  reg [31:0] _RAND_2200;
  reg [31:0] _RAND_2201;
  reg [31:0] _RAND_2202;
  reg [31:0] _RAND_2203;
  reg [31:0] _RAND_2204;
  reg [31:0] _RAND_2205;
  reg [31:0] _RAND_2206;
  reg [31:0] _RAND_2207;
  reg [31:0] _RAND_2208;
  reg [31:0] _RAND_2209;
  reg [31:0] _RAND_2210;
  reg [31:0] _RAND_2211;
  reg [31:0] _RAND_2212;
  reg [31:0] _RAND_2213;
  reg [31:0] _RAND_2214;
  reg [31:0] _RAND_2215;
  reg [31:0] _RAND_2216;
  reg [31:0] _RAND_2217;
  reg [31:0] _RAND_2218;
  reg [31:0] _RAND_2219;
  reg [31:0] _RAND_2220;
  reg [31:0] _RAND_2221;
  reg [31:0] _RAND_2222;
  reg [31:0] _RAND_2223;
  reg [31:0] _RAND_2224;
  reg [31:0] _RAND_2225;
  reg [31:0] _RAND_2226;
  reg [31:0] _RAND_2227;
  reg [31:0] _RAND_2228;
  reg [31:0] _RAND_2229;
  reg [31:0] _RAND_2230;
  reg [31:0] _RAND_2231;
  reg [31:0] _RAND_2232;
  reg [31:0] _RAND_2233;
  reg [31:0] _RAND_2234;
  reg [31:0] _RAND_2235;
  reg [31:0] _RAND_2236;
  reg [31:0] _RAND_2237;
  reg [31:0] _RAND_2238;
  reg [31:0] _RAND_2239;
  reg [31:0] _RAND_2240;
  reg [31:0] _RAND_2241;
  reg [31:0] _RAND_2242;
  reg [31:0] _RAND_2243;
  reg [31:0] _RAND_2244;
  reg [31:0] _RAND_2245;
  reg [31:0] _RAND_2246;
  reg [31:0] _RAND_2247;
  reg [31:0] _RAND_2248;
  reg [31:0] _RAND_2249;
  reg [31:0] _RAND_2250;
  reg [31:0] _RAND_2251;
  reg [31:0] _RAND_2252;
  reg [31:0] _RAND_2253;
  reg [31:0] _RAND_2254;
  reg [31:0] _RAND_2255;
  reg [31:0] _RAND_2256;
  reg [31:0] _RAND_2257;
  reg [31:0] _RAND_2258;
  reg [31:0] _RAND_2259;
  reg [31:0] _RAND_2260;
  reg [31:0] _RAND_2261;
  reg [31:0] _RAND_2262;
  reg [31:0] _RAND_2263;
  reg [31:0] _RAND_2264;
  reg [31:0] _RAND_2265;
  reg [31:0] _RAND_2266;
  reg [31:0] _RAND_2267;
  reg [31:0] _RAND_2268;
  reg [31:0] _RAND_2269;
  reg [31:0] _RAND_2270;
  reg [31:0] _RAND_2271;
  reg [31:0] _RAND_2272;
  reg [31:0] _RAND_2273;
  reg [31:0] _RAND_2274;
  reg [31:0] _RAND_2275;
  reg [31:0] _RAND_2276;
  reg [31:0] _RAND_2277;
  reg [31:0] _RAND_2278;
  reg [31:0] _RAND_2279;
  reg [31:0] _RAND_2280;
  reg [31:0] _RAND_2281;
  reg [31:0] _RAND_2282;
  reg [31:0] _RAND_2283;
  reg [31:0] _RAND_2284;
  reg [31:0] _RAND_2285;
  reg [31:0] _RAND_2286;
  reg [31:0] _RAND_2287;
  reg [31:0] _RAND_2288;
  reg [31:0] _RAND_2289;
  reg [31:0] _RAND_2290;
  reg [31:0] _RAND_2291;
  reg [31:0] _RAND_2292;
  reg [31:0] _RAND_2293;
  reg [31:0] _RAND_2294;
  reg [31:0] _RAND_2295;
  reg [31:0] _RAND_2296;
  reg [31:0] _RAND_2297;
  reg [31:0] _RAND_2298;
  reg [31:0] _RAND_2299;
  reg [31:0] _RAND_2300;
  reg [31:0] _RAND_2301;
  reg [31:0] _RAND_2302;
  reg [31:0] _RAND_2303;
  reg [31:0] _RAND_2304;
  reg [31:0] _RAND_2305;
  reg [31:0] _RAND_2306;
  reg [31:0] _RAND_2307;
  reg [31:0] _RAND_2308;
  reg [31:0] _RAND_2309;
  reg [31:0] _RAND_2310;
  reg [31:0] _RAND_2311;
  reg [31:0] _RAND_2312;
  reg [31:0] _RAND_2313;
  reg [31:0] _RAND_2314;
  reg [31:0] _RAND_2315;
  reg [31:0] _RAND_2316;
  reg [31:0] _RAND_2317;
  reg [31:0] _RAND_2318;
  reg [31:0] _RAND_2319;
  reg [31:0] _RAND_2320;
  reg [31:0] _RAND_2321;
  reg [31:0] _RAND_2322;
  reg [31:0] _RAND_2323;
  reg [31:0] _RAND_2324;
  reg [31:0] _RAND_2325;
  reg [31:0] _RAND_2326;
  reg [31:0] _RAND_2327;
  reg [31:0] _RAND_2328;
  reg [31:0] _RAND_2329;
  reg [31:0] _RAND_2330;
  reg [31:0] _RAND_2331;
  reg [31:0] _RAND_2332;
  reg [31:0] _RAND_2333;
  reg [31:0] _RAND_2334;
  reg [31:0] _RAND_2335;
  reg [31:0] _RAND_2336;
  reg [31:0] _RAND_2337;
  reg [31:0] _RAND_2338;
  reg [31:0] _RAND_2339;
  reg [31:0] _RAND_2340;
  reg [31:0] _RAND_2341;
  reg [31:0] _RAND_2342;
  reg [31:0] _RAND_2343;
  reg [31:0] _RAND_2344;
  reg [31:0] _RAND_2345;
  reg [31:0] _RAND_2346;
  reg [31:0] _RAND_2347;
  reg [31:0] _RAND_2348;
  reg [31:0] _RAND_2349;
  reg [31:0] _RAND_2350;
  reg [31:0] _RAND_2351;
  reg [31:0] _RAND_2352;
  reg [31:0] _RAND_2353;
  reg [31:0] _RAND_2354;
  reg [31:0] _RAND_2355;
  reg [31:0] _RAND_2356;
  reg [31:0] _RAND_2357;
  reg [31:0] _RAND_2358;
  reg [31:0] _RAND_2359;
  reg [31:0] _RAND_2360;
  reg [31:0] _RAND_2361;
  reg [31:0] _RAND_2362;
  reg [31:0] _RAND_2363;
  reg [31:0] _RAND_2364;
  reg [31:0] _RAND_2365;
  reg [31:0] _RAND_2366;
  reg [31:0] _RAND_2367;
  reg [31:0] _RAND_2368;
  reg [31:0] _RAND_2369;
  reg [31:0] _RAND_2370;
  reg [31:0] _RAND_2371;
  reg [31:0] _RAND_2372;
  reg [31:0] _RAND_2373;
  reg [31:0] _RAND_2374;
  reg [31:0] _RAND_2375;
  reg [31:0] _RAND_2376;
  reg [31:0] _RAND_2377;
  reg [31:0] _RAND_2378;
  reg [31:0] _RAND_2379;
  reg [31:0] _RAND_2380;
  reg [31:0] _RAND_2381;
  reg [31:0] _RAND_2382;
  reg [31:0] _RAND_2383;
  reg [31:0] _RAND_2384;
  reg [31:0] _RAND_2385;
  reg [31:0] _RAND_2386;
  reg [31:0] _RAND_2387;
  reg [31:0] _RAND_2388;
  reg [31:0] _RAND_2389;
  reg [31:0] _RAND_2390;
  reg [31:0] _RAND_2391;
  reg [31:0] _RAND_2392;
  reg [31:0] _RAND_2393;
  reg [31:0] _RAND_2394;
  reg [31:0] _RAND_2395;
  reg [31:0] _RAND_2396;
  reg [31:0] _RAND_2397;
  reg [31:0] _RAND_2398;
  reg [31:0] _RAND_2399;
  reg [31:0] _RAND_2400;
  reg [31:0] _RAND_2401;
  reg [31:0] _RAND_2402;
  reg [31:0] _RAND_2403;
  reg [31:0] _RAND_2404;
  reg [31:0] _RAND_2405;
  reg [31:0] _RAND_2406;
  reg [31:0] _RAND_2407;
  reg [31:0] _RAND_2408;
  reg [31:0] _RAND_2409;
  reg [31:0] _RAND_2410;
  reg [31:0] _RAND_2411;
  reg [31:0] _RAND_2412;
  reg [31:0] _RAND_2413;
  reg [31:0] _RAND_2414;
  reg [31:0] _RAND_2415;
  reg [31:0] _RAND_2416;
  reg [31:0] _RAND_2417;
  reg [31:0] _RAND_2418;
  reg [31:0] _RAND_2419;
  reg [31:0] _RAND_2420;
  reg [31:0] _RAND_2421;
  reg [31:0] _RAND_2422;
  reg [31:0] _RAND_2423;
  reg [31:0] _RAND_2424;
  reg [31:0] _RAND_2425;
  reg [31:0] _RAND_2426;
  reg [31:0] _RAND_2427;
  reg [31:0] _RAND_2428;
  reg [31:0] _RAND_2429;
  reg [31:0] _RAND_2430;
  reg [31:0] _RAND_2431;
  reg [31:0] _RAND_2432;
  reg [31:0] _RAND_2433;
  reg [31:0] _RAND_2434;
  reg [31:0] _RAND_2435;
  reg [31:0] _RAND_2436;
  reg [31:0] _RAND_2437;
  reg [31:0] _RAND_2438;
  reg [31:0] _RAND_2439;
  reg [31:0] _RAND_2440;
  reg [31:0] _RAND_2441;
  reg [31:0] _RAND_2442;
  reg [31:0] _RAND_2443;
  reg [31:0] _RAND_2444;
  reg [31:0] _RAND_2445;
  reg [31:0] _RAND_2446;
  reg [31:0] _RAND_2447;
  reg [31:0] _RAND_2448;
  reg [31:0] _RAND_2449;
  reg [31:0] _RAND_2450;
  reg [31:0] _RAND_2451;
  reg [31:0] _RAND_2452;
  reg [31:0] _RAND_2453;
  reg [31:0] _RAND_2454;
  reg [31:0] _RAND_2455;
  reg [31:0] _RAND_2456;
  reg [31:0] _RAND_2457;
  reg [31:0] _RAND_2458;
  reg [31:0] _RAND_2459;
  reg [31:0] _RAND_2460;
  reg [31:0] _RAND_2461;
  reg [31:0] _RAND_2462;
  reg [31:0] _RAND_2463;
  reg [31:0] _RAND_2464;
  reg [31:0] _RAND_2465;
  reg [31:0] _RAND_2466;
  reg [31:0] _RAND_2467;
  reg [31:0] _RAND_2468;
  reg [31:0] _RAND_2469;
  reg [31:0] _RAND_2470;
  reg [31:0] _RAND_2471;
  reg [31:0] _RAND_2472;
  reg [31:0] _RAND_2473;
  reg [31:0] _RAND_2474;
  reg [31:0] _RAND_2475;
  reg [31:0] _RAND_2476;
  reg [31:0] _RAND_2477;
  reg [31:0] _RAND_2478;
  reg [31:0] _RAND_2479;
  reg [31:0] _RAND_2480;
  reg [31:0] _RAND_2481;
  reg [31:0] _RAND_2482;
  reg [31:0] _RAND_2483;
  reg [31:0] _RAND_2484;
  reg [31:0] _RAND_2485;
  reg [31:0] _RAND_2486;
  reg [31:0] _RAND_2487;
  reg [31:0] _RAND_2488;
  reg [31:0] _RAND_2489;
  reg [31:0] _RAND_2490;
  reg [31:0] _RAND_2491;
  reg [31:0] _RAND_2492;
  reg [31:0] _RAND_2493;
  reg [31:0] _RAND_2494;
  reg [31:0] _RAND_2495;
  reg [31:0] _RAND_2496;
  reg [31:0] _RAND_2497;
  reg [31:0] _RAND_2498;
  reg [31:0] _RAND_2499;
  reg [31:0] _RAND_2500;
  reg [31:0] _RAND_2501;
  reg [31:0] _RAND_2502;
  reg [31:0] _RAND_2503;
  reg [31:0] _RAND_2504;
  reg [31:0] _RAND_2505;
  reg [31:0] _RAND_2506;
  reg [31:0] _RAND_2507;
  reg [31:0] _RAND_2508;
  reg [31:0] _RAND_2509;
  reg [31:0] _RAND_2510;
  reg [31:0] _RAND_2511;
  reg [31:0] _RAND_2512;
  reg [31:0] _RAND_2513;
  reg [31:0] _RAND_2514;
  reg [31:0] _RAND_2515;
  reg [31:0] _RAND_2516;
  reg [31:0] _RAND_2517;
  reg [31:0] _RAND_2518;
  reg [31:0] _RAND_2519;
  reg [31:0] _RAND_2520;
  reg [31:0] _RAND_2521;
  reg [31:0] _RAND_2522;
  reg [31:0] _RAND_2523;
  reg [31:0] _RAND_2524;
  reg [31:0] _RAND_2525;
  reg [31:0] _RAND_2526;
  reg [31:0] _RAND_2527;
  reg [31:0] _RAND_2528;
  reg [31:0] _RAND_2529;
  reg [31:0] _RAND_2530;
  reg [31:0] _RAND_2531;
  reg [31:0] _RAND_2532;
  reg [31:0] _RAND_2533;
  reg [31:0] _RAND_2534;
  reg [31:0] _RAND_2535;
  reg [31:0] _RAND_2536;
  reg [31:0] _RAND_2537;
  reg [31:0] _RAND_2538;
  reg [31:0] _RAND_2539;
  reg [31:0] _RAND_2540;
  reg [31:0] _RAND_2541;
  reg [31:0] _RAND_2542;
  reg [31:0] _RAND_2543;
  reg [31:0] _RAND_2544;
  reg [31:0] _RAND_2545;
  reg [31:0] _RAND_2546;
  reg [31:0] _RAND_2547;
  reg [31:0] _RAND_2548;
  reg [31:0] _RAND_2549;
  reg [31:0] _RAND_2550;
  reg [31:0] _RAND_2551;
  reg [31:0] _RAND_2552;
  reg [31:0] _RAND_2553;
  reg [31:0] _RAND_2554;
  reg [31:0] _RAND_2555;
  reg [31:0] _RAND_2556;
  reg [31:0] _RAND_2557;
  reg [31:0] _RAND_2558;
  reg [31:0] _RAND_2559;
  reg [31:0] _RAND_2560;
  reg [31:0] _RAND_2561;
  reg [31:0] _RAND_2562;
  reg [31:0] _RAND_2563;
  reg [31:0] _RAND_2564;
  reg [31:0] _RAND_2565;
  reg [31:0] _RAND_2566;
  reg [31:0] _RAND_2567;
  reg [31:0] _RAND_2568;
  reg [31:0] _RAND_2569;
  reg [31:0] _RAND_2570;
  reg [31:0] _RAND_2571;
  reg [31:0] _RAND_2572;
  reg [31:0] _RAND_2573;
  reg [31:0] _RAND_2574;
  reg [31:0] _RAND_2575;
  reg [31:0] _RAND_2576;
  reg [31:0] _RAND_2577;
  reg [31:0] _RAND_2578;
  reg [31:0] _RAND_2579;
  reg [31:0] _RAND_2580;
  reg [31:0] _RAND_2581;
  reg [31:0] _RAND_2582;
  reg [31:0] _RAND_2583;
  reg [31:0] _RAND_2584;
  reg [31:0] _RAND_2585;
  reg [31:0] _RAND_2586;
  reg [31:0] _RAND_2587;
  reg [31:0] _RAND_2588;
  reg [31:0] _RAND_2589;
  reg [31:0] _RAND_2590;
  reg [31:0] _RAND_2591;
  reg [31:0] _RAND_2592;
  reg [31:0] _RAND_2593;
  reg [31:0] _RAND_2594;
  reg [31:0] _RAND_2595;
  reg [31:0] _RAND_2596;
  reg [31:0] _RAND_2597;
  reg [31:0] _RAND_2598;
  reg [31:0] _RAND_2599;
  reg [31:0] _RAND_2600;
  reg [31:0] _RAND_2601;
  reg [31:0] _RAND_2602;
  reg [31:0] _RAND_2603;
  reg [31:0] _RAND_2604;
  reg [31:0] _RAND_2605;
  reg [31:0] _RAND_2606;
  reg [31:0] _RAND_2607;
  reg [31:0] _RAND_2608;
  reg [31:0] _RAND_2609;
  reg [31:0] _RAND_2610;
  reg [31:0] _RAND_2611;
  reg [31:0] _RAND_2612;
  reg [31:0] _RAND_2613;
  reg [31:0] _RAND_2614;
  reg [31:0] _RAND_2615;
  reg [31:0] _RAND_2616;
  reg [31:0] _RAND_2617;
  reg [31:0] _RAND_2618;
  reg [31:0] _RAND_2619;
  reg [31:0] _RAND_2620;
  reg [31:0] _RAND_2621;
  reg [31:0] _RAND_2622;
  reg [31:0] _RAND_2623;
  reg [31:0] _RAND_2624;
  reg [31:0] _RAND_2625;
  reg [31:0] _RAND_2626;
  reg [31:0] _RAND_2627;
  reg [31:0] _RAND_2628;
  reg [31:0] _RAND_2629;
  reg [31:0] _RAND_2630;
  reg [31:0] _RAND_2631;
  reg [31:0] _RAND_2632;
  reg [31:0] _RAND_2633;
  reg [31:0] _RAND_2634;
  reg [31:0] _RAND_2635;
  reg [31:0] _RAND_2636;
  reg [31:0] _RAND_2637;
  reg [31:0] _RAND_2638;
  reg [31:0] _RAND_2639;
  reg [31:0] _RAND_2640;
  reg [31:0] _RAND_2641;
  reg [31:0] _RAND_2642;
  reg [31:0] _RAND_2643;
  reg [31:0] _RAND_2644;
  reg [31:0] _RAND_2645;
  reg [31:0] _RAND_2646;
  reg [31:0] _RAND_2647;
  reg [31:0] _RAND_2648;
  reg [31:0] _RAND_2649;
  reg [31:0] _RAND_2650;
  reg [31:0] _RAND_2651;
  reg [31:0] _RAND_2652;
  reg [31:0] _RAND_2653;
  reg [31:0] _RAND_2654;
  reg [31:0] _RAND_2655;
  reg [31:0] _RAND_2656;
  reg [31:0] _RAND_2657;
  reg [31:0] _RAND_2658;
  reg [31:0] _RAND_2659;
  reg [31:0] _RAND_2660;
  reg [31:0] _RAND_2661;
  reg [31:0] _RAND_2662;
  reg [31:0] _RAND_2663;
  reg [31:0] _RAND_2664;
  reg [31:0] _RAND_2665;
  reg [31:0] _RAND_2666;
  reg [31:0] _RAND_2667;
  reg [31:0] _RAND_2668;
  reg [31:0] _RAND_2669;
  reg [31:0] _RAND_2670;
  reg [31:0] _RAND_2671;
  reg [31:0] _RAND_2672;
  reg [31:0] _RAND_2673;
  reg [31:0] _RAND_2674;
  reg [31:0] _RAND_2675;
  reg [31:0] _RAND_2676;
  reg [31:0] _RAND_2677;
  reg [31:0] _RAND_2678;
  reg [31:0] _RAND_2679;
  reg [31:0] _RAND_2680;
  reg [31:0] _RAND_2681;
  reg [31:0] _RAND_2682;
  reg [31:0] _RAND_2683;
  reg [31:0] _RAND_2684;
  reg [31:0] _RAND_2685;
  reg [31:0] _RAND_2686;
  reg [31:0] _RAND_2687;
  reg [31:0] _RAND_2688;
  reg [31:0] _RAND_2689;
  reg [31:0] _RAND_2690;
  reg [31:0] _RAND_2691;
  reg [31:0] _RAND_2692;
  reg [31:0] _RAND_2693;
  reg [31:0] _RAND_2694;
  reg [31:0] _RAND_2695;
  reg [31:0] _RAND_2696;
  reg [31:0] _RAND_2697;
  reg [31:0] _RAND_2698;
  reg [31:0] _RAND_2699;
  reg [31:0] _RAND_2700;
  reg [31:0] _RAND_2701;
  reg [31:0] _RAND_2702;
  reg [31:0] _RAND_2703;
  reg [31:0] _RAND_2704;
  reg [31:0] _RAND_2705;
  reg [31:0] _RAND_2706;
  reg [31:0] _RAND_2707;
  reg [31:0] _RAND_2708;
  reg [31:0] _RAND_2709;
  reg [31:0] _RAND_2710;
  reg [31:0] _RAND_2711;
  reg [31:0] _RAND_2712;
  reg [31:0] _RAND_2713;
  reg [31:0] _RAND_2714;
  reg [31:0] _RAND_2715;
  reg [31:0] _RAND_2716;
  reg [31:0] _RAND_2717;
  reg [31:0] _RAND_2718;
  reg [31:0] _RAND_2719;
  reg [31:0] _RAND_2720;
  reg [31:0] _RAND_2721;
  reg [31:0] _RAND_2722;
  reg [31:0] _RAND_2723;
  reg [31:0] _RAND_2724;
  reg [31:0] _RAND_2725;
  reg [31:0] _RAND_2726;
  reg [31:0] _RAND_2727;
  reg [31:0] _RAND_2728;
  reg [31:0] _RAND_2729;
  reg [31:0] _RAND_2730;
  reg [31:0] _RAND_2731;
  reg [31:0] _RAND_2732;
  reg [31:0] _RAND_2733;
  reg [31:0] _RAND_2734;
  reg [31:0] _RAND_2735;
  reg [31:0] _RAND_2736;
  reg [31:0] _RAND_2737;
  reg [31:0] _RAND_2738;
  reg [31:0] _RAND_2739;
  reg [31:0] _RAND_2740;
  reg [31:0] _RAND_2741;
  reg [31:0] _RAND_2742;
  reg [31:0] _RAND_2743;
  reg [31:0] _RAND_2744;
  reg [31:0] _RAND_2745;
  reg [31:0] _RAND_2746;
  reg [31:0] _RAND_2747;
  reg [31:0] _RAND_2748;
  reg [31:0] _RAND_2749;
  reg [31:0] _RAND_2750;
  reg [31:0] _RAND_2751;
  reg [31:0] _RAND_2752;
  reg [31:0] _RAND_2753;
  reg [31:0] _RAND_2754;
  reg [31:0] _RAND_2755;
  reg [31:0] _RAND_2756;
  reg [31:0] _RAND_2757;
  reg [31:0] _RAND_2758;
  reg [31:0] _RAND_2759;
  reg [31:0] _RAND_2760;
  reg [31:0] _RAND_2761;
  reg [31:0] _RAND_2762;
  reg [31:0] _RAND_2763;
  reg [31:0] _RAND_2764;
  reg [31:0] _RAND_2765;
  reg [31:0] _RAND_2766;
  reg [31:0] _RAND_2767;
  reg [31:0] _RAND_2768;
  reg [31:0] _RAND_2769;
  reg [31:0] _RAND_2770;
  reg [31:0] _RAND_2771;
  reg [31:0] _RAND_2772;
  reg [31:0] _RAND_2773;
  reg [31:0] _RAND_2774;
  reg [31:0] _RAND_2775;
  reg [31:0] _RAND_2776;
  reg [31:0] _RAND_2777;
  reg [31:0] _RAND_2778;
  reg [31:0] _RAND_2779;
  reg [31:0] _RAND_2780;
  reg [31:0] _RAND_2781;
  reg [31:0] _RAND_2782;
  reg [31:0] _RAND_2783;
  reg [31:0] _RAND_2784;
  reg [31:0] _RAND_2785;
  reg [31:0] _RAND_2786;
  reg [31:0] _RAND_2787;
  reg [31:0] _RAND_2788;
  reg [31:0] _RAND_2789;
  reg [31:0] _RAND_2790;
  reg [31:0] _RAND_2791;
  reg [31:0] _RAND_2792;
  reg [31:0] _RAND_2793;
  reg [31:0] _RAND_2794;
  reg [31:0] _RAND_2795;
  reg [31:0] _RAND_2796;
  reg [31:0] _RAND_2797;
  reg [31:0] _RAND_2798;
  reg [31:0] _RAND_2799;
  reg [31:0] _RAND_2800;
  reg [31:0] _RAND_2801;
  reg [31:0] _RAND_2802;
  reg [31:0] _RAND_2803;
  reg [31:0] _RAND_2804;
  reg [31:0] _RAND_2805;
  reg [31:0] _RAND_2806;
  reg [31:0] _RAND_2807;
  reg [31:0] _RAND_2808;
  reg [31:0] _RAND_2809;
  reg [31:0] _RAND_2810;
  reg [31:0] _RAND_2811;
  reg [31:0] _RAND_2812;
  reg [31:0] _RAND_2813;
  reg [31:0] _RAND_2814;
  reg [31:0] _RAND_2815;
  reg [31:0] _RAND_2816;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] Butterfly_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_1_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_1_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_1_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_1_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_1_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_2_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_2_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_2_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_2_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_2_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_3_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_3_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_3_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_3_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_3_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_4_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_4_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_4_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_4_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_4_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_5_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_5_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_5_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_5_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_5_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_6_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_6_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_6_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_6_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_6_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] Butterfly_7_io_in1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_in2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_wn_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out1_im; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_re; // @[Butterfly.scala 89:22]
  wire [31:0] Butterfly_7_io_out2_im; // @[Butterfly.scala 89:22]
  wire [31:0] Switch_7_io_in1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_in2_im; // @[Butterfly.scala 110:22]
  wire  Switch_7_io_sel; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out1_im; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_re; // @[Butterfly.scala 110:22]
  wire [31:0] Switch_7_io_out2_im; // @[Butterfly.scala 110:22]
  wire [31:0] ComplexAdd_io_op1_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op1_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_op2_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_re; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexAdd_io_res_im; // @[Butterfly.scala 26:22]
  wire [31:0] ComplexSub_io_op1_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op1_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_op2_im; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_re; // @[Butterfly.scala 40:22]
  wire [31:0] ComplexSub_io_res_im; // @[Butterfly.scala 40:22]
  reg [8:0] cnt; // @[FFT.scala 62:20]
  wire [8:0] _T_1 = cnt + 9'h1; // @[FFT.scala 64:16]
  wire [31:0] _GEN_2 = 8'h1 == cnt[7:0] ? $signed(32'shfffb) : $signed(32'sh10000); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3 = 8'h2 == cnt[7:0] ? $signed(32'shffec) : $signed(_GEN_2); // @[FFT.scala 51:18]
  wire [31:0] _GEN_4 = 8'h3 == cnt[7:0] ? $signed(32'shffd4) : $signed(_GEN_3); // @[FFT.scala 51:18]
  wire [31:0] _GEN_5 = 8'h4 == cnt[7:0] ? $signed(32'shffb1) : $signed(_GEN_4); // @[FFT.scala 51:18]
  wire [31:0] _GEN_6 = 8'h5 == cnt[7:0] ? $signed(32'shff85) : $signed(_GEN_5); // @[FFT.scala 51:18]
  wire [31:0] _GEN_7 = 8'h6 == cnt[7:0] ? $signed(32'shff4e) : $signed(_GEN_6); // @[FFT.scala 51:18]
  wire [31:0] _GEN_8 = 8'h7 == cnt[7:0] ? $signed(32'shff0e) : $signed(_GEN_7); // @[FFT.scala 51:18]
  wire [31:0] _GEN_9 = 8'h8 == cnt[7:0] ? $signed(32'shfec4) : $signed(_GEN_8); // @[FFT.scala 51:18]
  wire [31:0] _GEN_10 = 8'h9 == cnt[7:0] ? $signed(32'shfe71) : $signed(_GEN_9); // @[FFT.scala 51:18]
  wire [31:0] _GEN_11 = 8'ha == cnt[7:0] ? $signed(32'shfe13) : $signed(_GEN_10); // @[FFT.scala 51:18]
  wire [31:0] _GEN_12 = 8'hb == cnt[7:0] ? $signed(32'shfdac) : $signed(_GEN_11); // @[FFT.scala 51:18]
  wire [31:0] _GEN_13 = 8'hc == cnt[7:0] ? $signed(32'shfd3b) : $signed(_GEN_12); // @[FFT.scala 51:18]
  wire [31:0] _GEN_14 = 8'hd == cnt[7:0] ? $signed(32'shfcc0) : $signed(_GEN_13); // @[FFT.scala 51:18]
  wire [31:0] _GEN_15 = 8'he == cnt[7:0] ? $signed(32'shfc3b) : $signed(_GEN_14); // @[FFT.scala 51:18]
  wire [31:0] _GEN_16 = 8'hf == cnt[7:0] ? $signed(32'shfbad) : $signed(_GEN_15); // @[FFT.scala 51:18]
  wire [31:0] _GEN_17 = 8'h10 == cnt[7:0] ? $signed(32'shfb15) : $signed(_GEN_16); // @[FFT.scala 51:18]
  wire [31:0] _GEN_18 = 8'h11 == cnt[7:0] ? $signed(32'shfa73) : $signed(_GEN_17); // @[FFT.scala 51:18]
  wire [31:0] _GEN_19 = 8'h12 == cnt[7:0] ? $signed(32'shf9c8) : $signed(_GEN_18); // @[FFT.scala 51:18]
  wire [31:0] _GEN_20 = 8'h13 == cnt[7:0] ? $signed(32'shf913) : $signed(_GEN_19); // @[FFT.scala 51:18]
  wire [31:0] _GEN_21 = 8'h14 == cnt[7:0] ? $signed(32'shf854) : $signed(_GEN_20); // @[FFT.scala 51:18]
  wire [31:0] _GEN_22 = 8'h15 == cnt[7:0] ? $signed(32'shf78c) : $signed(_GEN_21); // @[FFT.scala 51:18]
  wire [31:0] _GEN_23 = 8'h16 == cnt[7:0] ? $signed(32'shf6ba) : $signed(_GEN_22); // @[FFT.scala 51:18]
  wire [31:0] _GEN_24 = 8'h17 == cnt[7:0] ? $signed(32'shf5df) : $signed(_GEN_23); // @[FFT.scala 51:18]
  wire [31:0] _GEN_25 = 8'h18 == cnt[7:0] ? $signed(32'shf4fa) : $signed(_GEN_24); // @[FFT.scala 51:18]
  wire [31:0] _GEN_26 = 8'h19 == cnt[7:0] ? $signed(32'shf40c) : $signed(_GEN_25); // @[FFT.scala 51:18]
  wire [31:0] _GEN_27 = 8'h1a == cnt[7:0] ? $signed(32'shf314) : $signed(_GEN_26); // @[FFT.scala 51:18]
  wire [31:0] _GEN_28 = 8'h1b == cnt[7:0] ? $signed(32'shf213) : $signed(_GEN_27); // @[FFT.scala 51:18]
  wire [31:0] _GEN_29 = 8'h1c == cnt[7:0] ? $signed(32'shf109) : $signed(_GEN_28); // @[FFT.scala 51:18]
  wire [31:0] _GEN_30 = 8'h1d == cnt[7:0] ? $signed(32'sheff5) : $signed(_GEN_29); // @[FFT.scala 51:18]
  wire [31:0] _GEN_31 = 8'h1e == cnt[7:0] ? $signed(32'sheed9) : $signed(_GEN_30); // @[FFT.scala 51:18]
  wire [31:0] _GEN_32 = 8'h1f == cnt[7:0] ? $signed(32'shedb3) : $signed(_GEN_31); // @[FFT.scala 51:18]
  wire [31:0] _GEN_33 = 8'h20 == cnt[7:0] ? $signed(32'shec83) : $signed(_GEN_32); // @[FFT.scala 51:18]
  wire [31:0] _GEN_34 = 8'h21 == cnt[7:0] ? $signed(32'sheb4b) : $signed(_GEN_33); // @[FFT.scala 51:18]
  wire [31:0] _GEN_35 = 8'h22 == cnt[7:0] ? $signed(32'shea0a) : $signed(_GEN_34); // @[FFT.scala 51:18]
  wire [31:0] _GEN_36 = 8'h23 == cnt[7:0] ? $signed(32'she8bf) : $signed(_GEN_35); // @[FFT.scala 51:18]
  wire [31:0] _GEN_37 = 8'h24 == cnt[7:0] ? $signed(32'she76c) : $signed(_GEN_36); // @[FFT.scala 51:18]
  wire [31:0] _GEN_38 = 8'h25 == cnt[7:0] ? $signed(32'she610) : $signed(_GEN_37); // @[FFT.scala 51:18]
  wire [31:0] _GEN_39 = 8'h26 == cnt[7:0] ? $signed(32'she4aa) : $signed(_GEN_38); // @[FFT.scala 51:18]
  wire [31:0] _GEN_40 = 8'h27 == cnt[7:0] ? $signed(32'she33c) : $signed(_GEN_39); // @[FFT.scala 51:18]
  wire [31:0] _GEN_41 = 8'h28 == cnt[7:0] ? $signed(32'she1c6) : $signed(_GEN_40); // @[FFT.scala 51:18]
  wire [31:0] _GEN_42 = 8'h29 == cnt[7:0] ? $signed(32'she046) : $signed(_GEN_41); // @[FFT.scala 51:18]
  wire [31:0] _GEN_43 = 8'h2a == cnt[7:0] ? $signed(32'shdebe) : $signed(_GEN_42); // @[FFT.scala 51:18]
  wire [31:0] _GEN_44 = 8'h2b == cnt[7:0] ? $signed(32'shdd2d) : $signed(_GEN_43); // @[FFT.scala 51:18]
  wire [31:0] _GEN_45 = 8'h2c == cnt[7:0] ? $signed(32'shdb94) : $signed(_GEN_44); // @[FFT.scala 51:18]
  wire [31:0] _GEN_46 = 8'h2d == cnt[7:0] ? $signed(32'shd9f2) : $signed(_GEN_45); // @[FFT.scala 51:18]
  wire [31:0] _GEN_47 = 8'h2e == cnt[7:0] ? $signed(32'shd848) : $signed(_GEN_46); // @[FFT.scala 51:18]
  wire [31:0] _GEN_48 = 8'h2f == cnt[7:0] ? $signed(32'shd696) : $signed(_GEN_47); // @[FFT.scala 51:18]
  wire [31:0] _GEN_49 = 8'h30 == cnt[7:0] ? $signed(32'shd4db) : $signed(_GEN_48); // @[FFT.scala 51:18]
  wire [31:0] _GEN_50 = 8'h31 == cnt[7:0] ? $signed(32'shd318) : $signed(_GEN_49); // @[FFT.scala 51:18]
  wire [31:0] _GEN_51 = 8'h32 == cnt[7:0] ? $signed(32'shd14d) : $signed(_GEN_50); // @[FFT.scala 51:18]
  wire [31:0] _GEN_52 = 8'h33 == cnt[7:0] ? $signed(32'shcf7a) : $signed(_GEN_51); // @[FFT.scala 51:18]
  wire [31:0] _GEN_53 = 8'h34 == cnt[7:0] ? $signed(32'shcd9f) : $signed(_GEN_52); // @[FFT.scala 51:18]
  wire [31:0] _GEN_54 = 8'h35 == cnt[7:0] ? $signed(32'shcbbc) : $signed(_GEN_53); // @[FFT.scala 51:18]
  wire [31:0] _GEN_55 = 8'h36 == cnt[7:0] ? $signed(32'shc9d1) : $signed(_GEN_54); // @[FFT.scala 51:18]
  wire [31:0] _GEN_56 = 8'h37 == cnt[7:0] ? $signed(32'shc7de) : $signed(_GEN_55); // @[FFT.scala 51:18]
  wire [31:0] _GEN_57 = 8'h38 == cnt[7:0] ? $signed(32'shc5e4) : $signed(_GEN_56); // @[FFT.scala 51:18]
  wire [31:0] _GEN_58 = 8'h39 == cnt[7:0] ? $signed(32'shc3e2) : $signed(_GEN_57); // @[FFT.scala 51:18]
  wire [31:0] _GEN_59 = 8'h3a == cnt[7:0] ? $signed(32'shc1d8) : $signed(_GEN_58); // @[FFT.scala 51:18]
  wire [31:0] _GEN_60 = 8'h3b == cnt[7:0] ? $signed(32'shbfc7) : $signed(_GEN_59); // @[FFT.scala 51:18]
  wire [31:0] _GEN_61 = 8'h3c == cnt[7:0] ? $signed(32'shbdaf) : $signed(_GEN_60); // @[FFT.scala 51:18]
  wire [31:0] _GEN_62 = 8'h3d == cnt[7:0] ? $signed(32'shbb8f) : $signed(_GEN_61); // @[FFT.scala 51:18]
  wire [31:0] _GEN_63 = 8'h3e == cnt[7:0] ? $signed(32'shb968) : $signed(_GEN_62); // @[FFT.scala 51:18]
  wire [31:0] _GEN_64 = 8'h3f == cnt[7:0] ? $signed(32'shb73a) : $signed(_GEN_63); // @[FFT.scala 51:18]
  wire [31:0] _GEN_65 = 8'h40 == cnt[7:0] ? $signed(32'shb505) : $signed(_GEN_64); // @[FFT.scala 51:18]
  wire [31:0] _GEN_66 = 8'h41 == cnt[7:0] ? $signed(32'shb2c9) : $signed(_GEN_65); // @[FFT.scala 51:18]
  wire [31:0] _GEN_67 = 8'h42 == cnt[7:0] ? $signed(32'shb086) : $signed(_GEN_66); // @[FFT.scala 51:18]
  wire [31:0] _GEN_68 = 8'h43 == cnt[7:0] ? $signed(32'shae3c) : $signed(_GEN_67); // @[FFT.scala 51:18]
  wire [31:0] _GEN_69 = 8'h44 == cnt[7:0] ? $signed(32'shabeb) : $signed(_GEN_68); // @[FFT.scala 51:18]
  wire [31:0] _GEN_70 = 8'h45 == cnt[7:0] ? $signed(32'sha994) : $signed(_GEN_69); // @[FFT.scala 51:18]
  wire [31:0] _GEN_71 = 8'h46 == cnt[7:0] ? $signed(32'sha736) : $signed(_GEN_70); // @[FFT.scala 51:18]
  wire [31:0] _GEN_72 = 8'h47 == cnt[7:0] ? $signed(32'sha4d2) : $signed(_GEN_71); // @[FFT.scala 51:18]
  wire [31:0] _GEN_73 = 8'h48 == cnt[7:0] ? $signed(32'sha268) : $signed(_GEN_72); // @[FFT.scala 51:18]
  wire [31:0] _GEN_74 = 8'h49 == cnt[7:0] ? $signed(32'sh9ff7) : $signed(_GEN_73); // @[FFT.scala 51:18]
  wire [31:0] _GEN_75 = 8'h4a == cnt[7:0] ? $signed(32'sh9d80) : $signed(_GEN_74); // @[FFT.scala 51:18]
  wire [31:0] _GEN_76 = 8'h4b == cnt[7:0] ? $signed(32'sh9b03) : $signed(_GEN_75); // @[FFT.scala 51:18]
  wire [31:0] _GEN_77 = 8'h4c == cnt[7:0] ? $signed(32'sh9880) : $signed(_GEN_76); // @[FFT.scala 51:18]
  wire [31:0] _GEN_78 = 8'h4d == cnt[7:0] ? $signed(32'sh95f7) : $signed(_GEN_77); // @[FFT.scala 51:18]
  wire [31:0] _GEN_79 = 8'h4e == cnt[7:0] ? $signed(32'sh9368) : $signed(_GEN_78); // @[FFT.scala 51:18]
  wire [31:0] _GEN_80 = 8'h4f == cnt[7:0] ? $signed(32'sh90d4) : $signed(_GEN_79); // @[FFT.scala 51:18]
  wire [31:0] _GEN_81 = 8'h50 == cnt[7:0] ? $signed(32'sh8e3a) : $signed(_GEN_80); // @[FFT.scala 51:18]
  wire [31:0] _GEN_82 = 8'h51 == cnt[7:0] ? $signed(32'sh8b9a) : $signed(_GEN_81); // @[FFT.scala 51:18]
  wire [31:0] _GEN_83 = 8'h52 == cnt[7:0] ? $signed(32'sh88f6) : $signed(_GEN_82); // @[FFT.scala 51:18]
  wire [31:0] _GEN_84 = 8'h53 == cnt[7:0] ? $signed(32'sh864c) : $signed(_GEN_83); // @[FFT.scala 51:18]
  wire [31:0] _GEN_85 = 8'h54 == cnt[7:0] ? $signed(32'sh839c) : $signed(_GEN_84); // @[FFT.scala 51:18]
  wire [31:0] _GEN_86 = 8'h55 == cnt[7:0] ? $signed(32'sh80e8) : $signed(_GEN_85); // @[FFT.scala 51:18]
  wire [31:0] _GEN_87 = 8'h56 == cnt[7:0] ? $signed(32'sh7e2f) : $signed(_GEN_86); // @[FFT.scala 51:18]
  wire [31:0] _GEN_88 = 8'h57 == cnt[7:0] ? $signed(32'sh7b70) : $signed(_GEN_87); // @[FFT.scala 51:18]
  wire [31:0] _GEN_89 = 8'h58 == cnt[7:0] ? $signed(32'sh78ad) : $signed(_GEN_88); // @[FFT.scala 51:18]
  wire [31:0] _GEN_90 = 8'h59 == cnt[7:0] ? $signed(32'sh75e6) : $signed(_GEN_89); // @[FFT.scala 51:18]
  wire [31:0] _GEN_91 = 8'h5a == cnt[7:0] ? $signed(32'sh731a) : $signed(_GEN_90); // @[FFT.scala 51:18]
  wire [31:0] _GEN_92 = 8'h5b == cnt[7:0] ? $signed(32'sh7049) : $signed(_GEN_91); // @[FFT.scala 51:18]
  wire [31:0] _GEN_93 = 8'h5c == cnt[7:0] ? $signed(32'sh6d74) : $signed(_GEN_92); // @[FFT.scala 51:18]
  wire [31:0] _GEN_94 = 8'h5d == cnt[7:0] ? $signed(32'sh6a9b) : $signed(_GEN_93); // @[FFT.scala 51:18]
  wire [31:0] _GEN_95 = 8'h5e == cnt[7:0] ? $signed(32'sh67be) : $signed(_GEN_94); // @[FFT.scala 51:18]
  wire [31:0] _GEN_96 = 8'h5f == cnt[7:0] ? $signed(32'sh64dd) : $signed(_GEN_95); // @[FFT.scala 51:18]
  wire [31:0] _GEN_97 = 8'h60 == cnt[7:0] ? $signed(32'sh61f8) : $signed(_GEN_96); // @[FFT.scala 51:18]
  wire [31:0] _GEN_98 = 8'h61 == cnt[7:0] ? $signed(32'sh5f0f) : $signed(_GEN_97); // @[FFT.scala 51:18]
  wire [31:0] _GEN_99 = 8'h62 == cnt[7:0] ? $signed(32'sh5c22) : $signed(_GEN_98); // @[FFT.scala 51:18]
  wire [31:0] _GEN_100 = 8'h63 == cnt[7:0] ? $signed(32'sh5932) : $signed(_GEN_99); // @[FFT.scala 51:18]
  wire [31:0] _GEN_101 = 8'h64 == cnt[7:0] ? $signed(32'sh563e) : $signed(_GEN_100); // @[FFT.scala 51:18]
  wire [31:0] _GEN_102 = 8'h65 == cnt[7:0] ? $signed(32'sh5348) : $signed(_GEN_101); // @[FFT.scala 51:18]
  wire [31:0] _GEN_103 = 8'h66 == cnt[7:0] ? $signed(32'sh504d) : $signed(_GEN_102); // @[FFT.scala 51:18]
  wire [31:0] _GEN_104 = 8'h67 == cnt[7:0] ? $signed(32'sh4d50) : $signed(_GEN_103); // @[FFT.scala 51:18]
  wire [31:0] _GEN_105 = 8'h68 == cnt[7:0] ? $signed(32'sh4a50) : $signed(_GEN_104); // @[FFT.scala 51:18]
  wire [31:0] _GEN_106 = 8'h69 == cnt[7:0] ? $signed(32'sh474d) : $signed(_GEN_105); // @[FFT.scala 51:18]
  wire [31:0] _GEN_107 = 8'h6a == cnt[7:0] ? $signed(32'sh4447) : $signed(_GEN_106); // @[FFT.scala 51:18]
  wire [31:0] _GEN_108 = 8'h6b == cnt[7:0] ? $signed(32'sh413f) : $signed(_GEN_107); // @[FFT.scala 51:18]
  wire [31:0] _GEN_109 = 8'h6c == cnt[7:0] ? $signed(32'sh3e34) : $signed(_GEN_108); // @[FFT.scala 51:18]
  wire [31:0] _GEN_110 = 8'h6d == cnt[7:0] ? $signed(32'sh3b27) : $signed(_GEN_109); // @[FFT.scala 51:18]
  wire [31:0] _GEN_111 = 8'h6e == cnt[7:0] ? $signed(32'sh3817) : $signed(_GEN_110); // @[FFT.scala 51:18]
  wire [31:0] _GEN_112 = 8'h6f == cnt[7:0] ? $signed(32'sh3505) : $signed(_GEN_111); // @[FFT.scala 51:18]
  wire [31:0] _GEN_113 = 8'h70 == cnt[7:0] ? $signed(32'sh31f1) : $signed(_GEN_112); // @[FFT.scala 51:18]
  wire [31:0] _GEN_114 = 8'h71 == cnt[7:0] ? $signed(32'sh2edc) : $signed(_GEN_113); // @[FFT.scala 51:18]
  wire [31:0] _GEN_115 = 8'h72 == cnt[7:0] ? $signed(32'sh2bc4) : $signed(_GEN_114); // @[FFT.scala 51:18]
  wire [31:0] _GEN_116 = 8'h73 == cnt[7:0] ? $signed(32'sh28ab) : $signed(_GEN_115); // @[FFT.scala 51:18]
  wire [31:0] _GEN_117 = 8'h74 == cnt[7:0] ? $signed(32'sh2590) : $signed(_GEN_116); // @[FFT.scala 51:18]
  wire [31:0] _GEN_118 = 8'h75 == cnt[7:0] ? $signed(32'sh2274) : $signed(_GEN_117); // @[FFT.scala 51:18]
  wire [31:0] _GEN_119 = 8'h76 == cnt[7:0] ? $signed(32'sh1f56) : $signed(_GEN_118); // @[FFT.scala 51:18]
  wire [31:0] _GEN_120 = 8'h77 == cnt[7:0] ? $signed(32'sh1c38) : $signed(_GEN_119); // @[FFT.scala 51:18]
  wire [31:0] _GEN_121 = 8'h78 == cnt[7:0] ? $signed(32'sh1918) : $signed(_GEN_120); // @[FFT.scala 51:18]
  wire [31:0] _GEN_122 = 8'h79 == cnt[7:0] ? $signed(32'sh15f7) : $signed(_GEN_121); // @[FFT.scala 51:18]
  wire [31:0] _GEN_123 = 8'h7a == cnt[7:0] ? $signed(32'sh12d5) : $signed(_GEN_122); // @[FFT.scala 51:18]
  wire [31:0] _GEN_124 = 8'h7b == cnt[7:0] ? $signed(32'shfb3) : $signed(_GEN_123); // @[FFT.scala 51:18]
  wire [31:0] _GEN_125 = 8'h7c == cnt[7:0] ? $signed(32'shc90) : $signed(_GEN_124); // @[FFT.scala 51:18]
  wire [31:0] _GEN_126 = 8'h7d == cnt[7:0] ? $signed(32'sh96c) : $signed(_GEN_125); // @[FFT.scala 51:18]
  wire [31:0] _GEN_127 = 8'h7e == cnt[7:0] ? $signed(32'sh648) : $signed(_GEN_126); // @[FFT.scala 51:18]
  wire [31:0] _GEN_128 = 8'h7f == cnt[7:0] ? $signed(32'sh324) : $signed(_GEN_127); // @[FFT.scala 51:18]
  wire [31:0] _GEN_129 = 8'h80 == cnt[7:0] ? $signed(32'sh0) : $signed(_GEN_128); // @[FFT.scala 51:18]
  wire [31:0] _GEN_130 = 8'h81 == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_129); // @[FFT.scala 51:18]
  wire [31:0] _GEN_131 = 8'h82 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_130); // @[FFT.scala 51:18]
  wire [31:0] _GEN_132 = 8'h83 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_131); // @[FFT.scala 51:18]
  wire [31:0] _GEN_133 = 8'h84 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_132); // @[FFT.scala 51:18]
  wire [31:0] _GEN_134 = 8'h85 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_133); // @[FFT.scala 51:18]
  wire [31:0] _GEN_135 = 8'h86 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_134); // @[FFT.scala 51:18]
  wire [31:0] _GEN_136 = 8'h87 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_135); // @[FFT.scala 51:18]
  wire [31:0] _GEN_137 = 8'h88 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_136); // @[FFT.scala 51:18]
  wire [31:0] _GEN_138 = 8'h89 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_137); // @[FFT.scala 51:18]
  wire [31:0] _GEN_139 = 8'h8a == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_138); // @[FFT.scala 51:18]
  wire [31:0] _GEN_140 = 8'h8b == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_139); // @[FFT.scala 51:18]
  wire [31:0] _GEN_141 = 8'h8c == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_140); // @[FFT.scala 51:18]
  wire [31:0] _GEN_142 = 8'h8d == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_141); // @[FFT.scala 51:18]
  wire [31:0] _GEN_143 = 8'h8e == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_142); // @[FFT.scala 51:18]
  wire [31:0] _GEN_144 = 8'h8f == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_143); // @[FFT.scala 51:18]
  wire [31:0] _GEN_145 = 8'h90 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_144); // @[FFT.scala 51:18]
  wire [31:0] _GEN_146 = 8'h91 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_145); // @[FFT.scala 51:18]
  wire [31:0] _GEN_147 = 8'h92 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_146); // @[FFT.scala 51:18]
  wire [31:0] _GEN_148 = 8'h93 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_147); // @[FFT.scala 51:18]
  wire [31:0] _GEN_149 = 8'h94 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_148); // @[FFT.scala 51:18]
  wire [31:0] _GEN_150 = 8'h95 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_149); // @[FFT.scala 51:18]
  wire [31:0] _GEN_151 = 8'h96 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_150); // @[FFT.scala 51:18]
  wire [31:0] _GEN_152 = 8'h97 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_151); // @[FFT.scala 51:18]
  wire [31:0] _GEN_153 = 8'h98 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_152); // @[FFT.scala 51:18]
  wire [31:0] _GEN_154 = 8'h99 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_153); // @[FFT.scala 51:18]
  wire [31:0] _GEN_155 = 8'h9a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_154); // @[FFT.scala 51:18]
  wire [31:0] _GEN_156 = 8'h9b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_155); // @[FFT.scala 51:18]
  wire [31:0] _GEN_157 = 8'h9c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_156); // @[FFT.scala 51:18]
  wire [31:0] _GEN_158 = 8'h9d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_157); // @[FFT.scala 51:18]
  wire [31:0] _GEN_159 = 8'h9e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_158); // @[FFT.scala 51:18]
  wire [31:0] _GEN_160 = 8'h9f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_159); // @[FFT.scala 51:18]
  wire [31:0] _GEN_161 = 8'ha0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_160); // @[FFT.scala 51:18]
  wire [31:0] _GEN_162 = 8'ha1 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_161); // @[FFT.scala 51:18]
  wire [31:0] _GEN_163 = 8'ha2 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_162); // @[FFT.scala 51:18]
  wire [31:0] _GEN_164 = 8'ha3 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_163); // @[FFT.scala 51:18]
  wire [31:0] _GEN_165 = 8'ha4 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_164); // @[FFT.scala 51:18]
  wire [31:0] _GEN_166 = 8'ha5 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_165); // @[FFT.scala 51:18]
  wire [31:0] _GEN_167 = 8'ha6 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_166); // @[FFT.scala 51:18]
  wire [31:0] _GEN_168 = 8'ha7 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_167); // @[FFT.scala 51:18]
  wire [31:0] _GEN_169 = 8'ha8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_168); // @[FFT.scala 51:18]
  wire [31:0] _GEN_170 = 8'ha9 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_169); // @[FFT.scala 51:18]
  wire [31:0] _GEN_171 = 8'haa == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_170); // @[FFT.scala 51:18]
  wire [31:0] _GEN_172 = 8'hab == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_171); // @[FFT.scala 51:18]
  wire [31:0] _GEN_173 = 8'hac == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_172); // @[FFT.scala 51:18]
  wire [31:0] _GEN_174 = 8'had == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_173); // @[FFT.scala 51:18]
  wire [31:0] _GEN_175 = 8'hae == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_174); // @[FFT.scala 51:18]
  wire [31:0] _GEN_176 = 8'haf == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_175); // @[FFT.scala 51:18]
  wire [31:0] _GEN_177 = 8'hb0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_176); // @[FFT.scala 51:18]
  wire [31:0] _GEN_178 = 8'hb1 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_177); // @[FFT.scala 51:18]
  wire [31:0] _GEN_179 = 8'hb2 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_178); // @[FFT.scala 51:18]
  wire [31:0] _GEN_180 = 8'hb3 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_179); // @[FFT.scala 51:18]
  wire [31:0] _GEN_181 = 8'hb4 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_180); // @[FFT.scala 51:18]
  wire [31:0] _GEN_182 = 8'hb5 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_181); // @[FFT.scala 51:18]
  wire [31:0] _GEN_183 = 8'hb6 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_182); // @[FFT.scala 51:18]
  wire [31:0] _GEN_184 = 8'hb7 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_183); // @[FFT.scala 51:18]
  wire [31:0] _GEN_185 = 8'hb8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_184); // @[FFT.scala 51:18]
  wire [31:0] _GEN_186 = 8'hb9 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_185); // @[FFT.scala 51:18]
  wire [31:0] _GEN_187 = 8'hba == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_186); // @[FFT.scala 51:18]
  wire [31:0] _GEN_188 = 8'hbb == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_187); // @[FFT.scala 51:18]
  wire [31:0] _GEN_189 = 8'hbc == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_188); // @[FFT.scala 51:18]
  wire [31:0] _GEN_190 = 8'hbd == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_189); // @[FFT.scala 51:18]
  wire [31:0] _GEN_191 = 8'hbe == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_190); // @[FFT.scala 51:18]
  wire [31:0] _GEN_192 = 8'hbf == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_191); // @[FFT.scala 51:18]
  wire [31:0] _GEN_193 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_192); // @[FFT.scala 51:18]
  wire [31:0] _GEN_194 = 8'hc1 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_193); // @[FFT.scala 51:18]
  wire [31:0] _GEN_195 = 8'hc2 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_194); // @[FFT.scala 51:18]
  wire [31:0] _GEN_196 = 8'hc3 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_195); // @[FFT.scala 51:18]
  wire [31:0] _GEN_197 = 8'hc4 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_196); // @[FFT.scala 51:18]
  wire [31:0] _GEN_198 = 8'hc5 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_197); // @[FFT.scala 51:18]
  wire [31:0] _GEN_199 = 8'hc6 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_198); // @[FFT.scala 51:18]
  wire [31:0] _GEN_200 = 8'hc7 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_199); // @[FFT.scala 51:18]
  wire [31:0] _GEN_201 = 8'hc8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_200); // @[FFT.scala 51:18]
  wire [31:0] _GEN_202 = 8'hc9 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_201); // @[FFT.scala 51:18]
  wire [31:0] _GEN_203 = 8'hca == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_202); // @[FFT.scala 51:18]
  wire [31:0] _GEN_204 = 8'hcb == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_203); // @[FFT.scala 51:18]
  wire [31:0] _GEN_205 = 8'hcc == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_204); // @[FFT.scala 51:18]
  wire [31:0] _GEN_206 = 8'hcd == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_205); // @[FFT.scala 51:18]
  wire [31:0] _GEN_207 = 8'hce == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_206); // @[FFT.scala 51:18]
  wire [31:0] _GEN_208 = 8'hcf == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_207); // @[FFT.scala 51:18]
  wire [31:0] _GEN_209 = 8'hd0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_208); // @[FFT.scala 51:18]
  wire [31:0] _GEN_210 = 8'hd1 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_209); // @[FFT.scala 51:18]
  wire [31:0] _GEN_211 = 8'hd2 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_210); // @[FFT.scala 51:18]
  wire [31:0] _GEN_212 = 8'hd3 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_211); // @[FFT.scala 51:18]
  wire [31:0] _GEN_213 = 8'hd4 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_212); // @[FFT.scala 51:18]
  wire [31:0] _GEN_214 = 8'hd5 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_213); // @[FFT.scala 51:18]
  wire [31:0] _GEN_215 = 8'hd6 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_214); // @[FFT.scala 51:18]
  wire [31:0] _GEN_216 = 8'hd7 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_215); // @[FFT.scala 51:18]
  wire [31:0] _GEN_217 = 8'hd8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_216); // @[FFT.scala 51:18]
  wire [31:0] _GEN_218 = 8'hd9 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_217); // @[FFT.scala 51:18]
  wire [31:0] _GEN_219 = 8'hda == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_218); // @[FFT.scala 51:18]
  wire [31:0] _GEN_220 = 8'hdb == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_219); // @[FFT.scala 51:18]
  wire [31:0] _GEN_221 = 8'hdc == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_220); // @[FFT.scala 51:18]
  wire [31:0] _GEN_222 = 8'hdd == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_221); // @[FFT.scala 51:18]
  wire [31:0] _GEN_223 = 8'hde == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_222); // @[FFT.scala 51:18]
  wire [31:0] _GEN_224 = 8'hdf == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_223); // @[FFT.scala 51:18]
  wire [31:0] _GEN_225 = 8'he0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_224); // @[FFT.scala 51:18]
  wire [31:0] _GEN_226 = 8'he1 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_225); // @[FFT.scala 51:18]
  wire [31:0] _GEN_227 = 8'he2 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_226); // @[FFT.scala 51:18]
  wire [31:0] _GEN_228 = 8'he3 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_227); // @[FFT.scala 51:18]
  wire [31:0] _GEN_229 = 8'he4 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_228); // @[FFT.scala 51:18]
  wire [31:0] _GEN_230 = 8'he5 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_229); // @[FFT.scala 51:18]
  wire [31:0] _GEN_231 = 8'he6 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_230); // @[FFT.scala 51:18]
  wire [31:0] _GEN_232 = 8'he7 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_231); // @[FFT.scala 51:18]
  wire [31:0] _GEN_233 = 8'he8 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_232); // @[FFT.scala 51:18]
  wire [31:0] _GEN_234 = 8'he9 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_233); // @[FFT.scala 51:18]
  wire [31:0] _GEN_235 = 8'hea == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_234); // @[FFT.scala 51:18]
  wire [31:0] _GEN_236 = 8'heb == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_235); // @[FFT.scala 51:18]
  wire [31:0] _GEN_237 = 8'hec == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_236); // @[FFT.scala 51:18]
  wire [31:0] _GEN_238 = 8'hed == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_237); // @[FFT.scala 51:18]
  wire [31:0] _GEN_239 = 8'hee == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_238); // @[FFT.scala 51:18]
  wire [31:0] _GEN_240 = 8'hef == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_239); // @[FFT.scala 51:18]
  wire [31:0] _GEN_241 = 8'hf0 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_240); // @[FFT.scala 51:18]
  wire [31:0] _GEN_242 = 8'hf1 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_241); // @[FFT.scala 51:18]
  wire [31:0] _GEN_243 = 8'hf2 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_242); // @[FFT.scala 51:18]
  wire [31:0] _GEN_244 = 8'hf3 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_243); // @[FFT.scala 51:18]
  wire [31:0] _GEN_245 = 8'hf4 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_244); // @[FFT.scala 51:18]
  wire [31:0] _GEN_246 = 8'hf5 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_245); // @[FFT.scala 51:18]
  wire [31:0] _GEN_247 = 8'hf6 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_246); // @[FFT.scala 51:18]
  wire [31:0] _GEN_248 = 8'hf7 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_247); // @[FFT.scala 51:18]
  wire [31:0] _GEN_249 = 8'hf8 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_248); // @[FFT.scala 51:18]
  wire [31:0] _GEN_250 = 8'hf9 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_249); // @[FFT.scala 51:18]
  wire [31:0] _GEN_251 = 8'hfa == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_250); // @[FFT.scala 51:18]
  wire [31:0] _GEN_252 = 8'hfb == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_251); // @[FFT.scala 51:18]
  wire [31:0] _GEN_253 = 8'hfc == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_252); // @[FFT.scala 51:18]
  wire [31:0] _GEN_254 = 8'hfd == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_253); // @[FFT.scala 51:18]
  wire [31:0] _GEN_255 = 8'hfe == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_254); // @[FFT.scala 51:18]
  wire [31:0] _GEN_770 = 8'h1 == cnt[7:0] ? $signed(-32'sh324) : $signed(32'sh0); // @[FFT.scala 52:18]
  wire [31:0] _GEN_771 = 8'h2 == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_770); // @[FFT.scala 52:18]
  wire [31:0] _GEN_772 = 8'h3 == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_771); // @[FFT.scala 52:18]
  wire [31:0] _GEN_773 = 8'h4 == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_772); // @[FFT.scala 52:18]
  wire [31:0] _GEN_774 = 8'h5 == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_773); // @[FFT.scala 52:18]
  wire [31:0] _GEN_775 = 8'h6 == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_774); // @[FFT.scala 52:18]
  wire [31:0] _GEN_776 = 8'h7 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_775); // @[FFT.scala 52:18]
  wire [31:0] _GEN_777 = 8'h8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_776); // @[FFT.scala 52:18]
  wire [31:0] _GEN_778 = 8'h9 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_777); // @[FFT.scala 52:18]
  wire [31:0] _GEN_779 = 8'ha == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_778); // @[FFT.scala 52:18]
  wire [31:0] _GEN_780 = 8'hb == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_779); // @[FFT.scala 52:18]
  wire [31:0] _GEN_781 = 8'hc == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_780); // @[FFT.scala 52:18]
  wire [31:0] _GEN_782 = 8'hd == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_781); // @[FFT.scala 52:18]
  wire [31:0] _GEN_783 = 8'he == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_782); // @[FFT.scala 52:18]
  wire [31:0] _GEN_784 = 8'hf == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_783); // @[FFT.scala 52:18]
  wire [31:0] _GEN_785 = 8'h10 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_784); // @[FFT.scala 52:18]
  wire [31:0] _GEN_786 = 8'h11 == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_785); // @[FFT.scala 52:18]
  wire [31:0] _GEN_787 = 8'h12 == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_786); // @[FFT.scala 52:18]
  wire [31:0] _GEN_788 = 8'h13 == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_787); // @[FFT.scala 52:18]
  wire [31:0] _GEN_789 = 8'h14 == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_788); // @[FFT.scala 52:18]
  wire [31:0] _GEN_790 = 8'h15 == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_789); // @[FFT.scala 52:18]
  wire [31:0] _GEN_791 = 8'h16 == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_790); // @[FFT.scala 52:18]
  wire [31:0] _GEN_792 = 8'h17 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_791); // @[FFT.scala 52:18]
  wire [31:0] _GEN_793 = 8'h18 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_792); // @[FFT.scala 52:18]
  wire [31:0] _GEN_794 = 8'h19 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_793); // @[FFT.scala 52:18]
  wire [31:0] _GEN_795 = 8'h1a == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_794); // @[FFT.scala 52:18]
  wire [31:0] _GEN_796 = 8'h1b == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_795); // @[FFT.scala 52:18]
  wire [31:0] _GEN_797 = 8'h1c == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_796); // @[FFT.scala 52:18]
  wire [31:0] _GEN_798 = 8'h1d == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_797); // @[FFT.scala 52:18]
  wire [31:0] _GEN_799 = 8'h1e == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_798); // @[FFT.scala 52:18]
  wire [31:0] _GEN_800 = 8'h1f == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_799); // @[FFT.scala 52:18]
  wire [31:0] _GEN_801 = 8'h20 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_800); // @[FFT.scala 52:18]
  wire [31:0] _GEN_802 = 8'h21 == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_801); // @[FFT.scala 52:18]
  wire [31:0] _GEN_803 = 8'h22 == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_802); // @[FFT.scala 52:18]
  wire [31:0] _GEN_804 = 8'h23 == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_803); // @[FFT.scala 52:18]
  wire [31:0] _GEN_805 = 8'h24 == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_804); // @[FFT.scala 52:18]
  wire [31:0] _GEN_806 = 8'h25 == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_805); // @[FFT.scala 52:18]
  wire [31:0] _GEN_807 = 8'h26 == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_806); // @[FFT.scala 52:18]
  wire [31:0] _GEN_808 = 8'h27 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_807); // @[FFT.scala 52:18]
  wire [31:0] _GEN_809 = 8'h28 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_808); // @[FFT.scala 52:18]
  wire [31:0] _GEN_810 = 8'h29 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_809); // @[FFT.scala 52:18]
  wire [31:0] _GEN_811 = 8'h2a == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_810); // @[FFT.scala 52:18]
  wire [31:0] _GEN_812 = 8'h2b == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_811); // @[FFT.scala 52:18]
  wire [31:0] _GEN_813 = 8'h2c == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_812); // @[FFT.scala 52:18]
  wire [31:0] _GEN_814 = 8'h2d == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_813); // @[FFT.scala 52:18]
  wire [31:0] _GEN_815 = 8'h2e == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_814); // @[FFT.scala 52:18]
  wire [31:0] _GEN_816 = 8'h2f == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_815); // @[FFT.scala 52:18]
  wire [31:0] _GEN_817 = 8'h30 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_816); // @[FFT.scala 52:18]
  wire [31:0] _GEN_818 = 8'h31 == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_817); // @[FFT.scala 52:18]
  wire [31:0] _GEN_819 = 8'h32 == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_818); // @[FFT.scala 52:18]
  wire [31:0] _GEN_820 = 8'h33 == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_819); // @[FFT.scala 52:18]
  wire [31:0] _GEN_821 = 8'h34 == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_820); // @[FFT.scala 52:18]
  wire [31:0] _GEN_822 = 8'h35 == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_821); // @[FFT.scala 52:18]
  wire [31:0] _GEN_823 = 8'h36 == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_822); // @[FFT.scala 52:18]
  wire [31:0] _GEN_824 = 8'h37 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_823); // @[FFT.scala 52:18]
  wire [31:0] _GEN_825 = 8'h38 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_824); // @[FFT.scala 52:18]
  wire [31:0] _GEN_826 = 8'h39 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_825); // @[FFT.scala 52:18]
  wire [31:0] _GEN_827 = 8'h3a == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_826); // @[FFT.scala 52:18]
  wire [31:0] _GEN_828 = 8'h3b == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_827); // @[FFT.scala 52:18]
  wire [31:0] _GEN_829 = 8'h3c == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_828); // @[FFT.scala 52:18]
  wire [31:0] _GEN_830 = 8'h3d == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_829); // @[FFT.scala 52:18]
  wire [31:0] _GEN_831 = 8'h3e == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_830); // @[FFT.scala 52:18]
  wire [31:0] _GEN_832 = 8'h3f == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_831); // @[FFT.scala 52:18]
  wire [31:0] _GEN_833 = 8'h40 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_832); // @[FFT.scala 52:18]
  wire [31:0] _GEN_834 = 8'h41 == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_833); // @[FFT.scala 52:18]
  wire [31:0] _GEN_835 = 8'h42 == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_834); // @[FFT.scala 52:18]
  wire [31:0] _GEN_836 = 8'h43 == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_835); // @[FFT.scala 52:18]
  wire [31:0] _GEN_837 = 8'h44 == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_836); // @[FFT.scala 52:18]
  wire [31:0] _GEN_838 = 8'h45 == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_837); // @[FFT.scala 52:18]
  wire [31:0] _GEN_839 = 8'h46 == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_838); // @[FFT.scala 52:18]
  wire [31:0] _GEN_840 = 8'h47 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_839); // @[FFT.scala 52:18]
  wire [31:0] _GEN_841 = 8'h48 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_840); // @[FFT.scala 52:18]
  wire [31:0] _GEN_842 = 8'h49 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_841); // @[FFT.scala 52:18]
  wire [31:0] _GEN_843 = 8'h4a == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_842); // @[FFT.scala 52:18]
  wire [31:0] _GEN_844 = 8'h4b == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_843); // @[FFT.scala 52:18]
  wire [31:0] _GEN_845 = 8'h4c == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_844); // @[FFT.scala 52:18]
  wire [31:0] _GEN_846 = 8'h4d == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_845); // @[FFT.scala 52:18]
  wire [31:0] _GEN_847 = 8'h4e == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_846); // @[FFT.scala 52:18]
  wire [31:0] _GEN_848 = 8'h4f == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_847); // @[FFT.scala 52:18]
  wire [31:0] _GEN_849 = 8'h50 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_848); // @[FFT.scala 52:18]
  wire [31:0] _GEN_850 = 8'h51 == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_849); // @[FFT.scala 52:18]
  wire [31:0] _GEN_851 = 8'h52 == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_850); // @[FFT.scala 52:18]
  wire [31:0] _GEN_852 = 8'h53 == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_851); // @[FFT.scala 52:18]
  wire [31:0] _GEN_853 = 8'h54 == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_852); // @[FFT.scala 52:18]
  wire [31:0] _GEN_854 = 8'h55 == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_853); // @[FFT.scala 52:18]
  wire [31:0] _GEN_855 = 8'h56 == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_854); // @[FFT.scala 52:18]
  wire [31:0] _GEN_856 = 8'h57 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_855); // @[FFT.scala 52:18]
  wire [31:0] _GEN_857 = 8'h58 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_856); // @[FFT.scala 52:18]
  wire [31:0] _GEN_858 = 8'h59 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_857); // @[FFT.scala 52:18]
  wire [31:0] _GEN_859 = 8'h5a == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_858); // @[FFT.scala 52:18]
  wire [31:0] _GEN_860 = 8'h5b == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_859); // @[FFT.scala 52:18]
  wire [31:0] _GEN_861 = 8'h5c == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_860); // @[FFT.scala 52:18]
  wire [31:0] _GEN_862 = 8'h5d == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_861); // @[FFT.scala 52:18]
  wire [31:0] _GEN_863 = 8'h5e == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_862); // @[FFT.scala 52:18]
  wire [31:0] _GEN_864 = 8'h5f == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_863); // @[FFT.scala 52:18]
  wire [31:0] _GEN_865 = 8'h60 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_864); // @[FFT.scala 52:18]
  wire [31:0] _GEN_866 = 8'h61 == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_865); // @[FFT.scala 52:18]
  wire [31:0] _GEN_867 = 8'h62 == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_866); // @[FFT.scala 52:18]
  wire [31:0] _GEN_868 = 8'h63 == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_867); // @[FFT.scala 52:18]
  wire [31:0] _GEN_869 = 8'h64 == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_868); // @[FFT.scala 52:18]
  wire [31:0] _GEN_870 = 8'h65 == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_869); // @[FFT.scala 52:18]
  wire [31:0] _GEN_871 = 8'h66 == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_870); // @[FFT.scala 52:18]
  wire [31:0] _GEN_872 = 8'h67 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_871); // @[FFT.scala 52:18]
  wire [31:0] _GEN_873 = 8'h68 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_872); // @[FFT.scala 52:18]
  wire [31:0] _GEN_874 = 8'h69 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_873); // @[FFT.scala 52:18]
  wire [31:0] _GEN_875 = 8'h6a == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_874); // @[FFT.scala 52:18]
  wire [31:0] _GEN_876 = 8'h6b == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_875); // @[FFT.scala 52:18]
  wire [31:0] _GEN_877 = 8'h6c == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_876); // @[FFT.scala 52:18]
  wire [31:0] _GEN_878 = 8'h6d == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_877); // @[FFT.scala 52:18]
  wire [31:0] _GEN_879 = 8'h6e == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_878); // @[FFT.scala 52:18]
  wire [31:0] _GEN_880 = 8'h6f == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_879); // @[FFT.scala 52:18]
  wire [31:0] _GEN_881 = 8'h70 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_880); // @[FFT.scala 52:18]
  wire [31:0] _GEN_882 = 8'h71 == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_881); // @[FFT.scala 52:18]
  wire [31:0] _GEN_883 = 8'h72 == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_882); // @[FFT.scala 52:18]
  wire [31:0] _GEN_884 = 8'h73 == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_883); // @[FFT.scala 52:18]
  wire [31:0] _GEN_885 = 8'h74 == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_884); // @[FFT.scala 52:18]
  wire [31:0] _GEN_886 = 8'h75 == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_885); // @[FFT.scala 52:18]
  wire [31:0] _GEN_887 = 8'h76 == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_886); // @[FFT.scala 52:18]
  wire [31:0] _GEN_888 = 8'h77 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_887); // @[FFT.scala 52:18]
  wire [31:0] _GEN_889 = 8'h78 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_888); // @[FFT.scala 52:18]
  wire [31:0] _GEN_890 = 8'h79 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_889); // @[FFT.scala 52:18]
  wire [31:0] _GEN_891 = 8'h7a == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_890); // @[FFT.scala 52:18]
  wire [31:0] _GEN_892 = 8'h7b == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_891); // @[FFT.scala 52:18]
  wire [31:0] _GEN_893 = 8'h7c == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_892); // @[FFT.scala 52:18]
  wire [31:0] _GEN_894 = 8'h7d == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_893); // @[FFT.scala 52:18]
  wire [31:0] _GEN_895 = 8'h7e == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_894); // @[FFT.scala 52:18]
  wire [31:0] _GEN_896 = 8'h7f == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_895); // @[FFT.scala 52:18]
  wire [31:0] _GEN_897 = 8'h80 == cnt[7:0] ? $signed(-32'sh10000) : $signed(_GEN_896); // @[FFT.scala 52:18]
  wire [31:0] _GEN_898 = 8'h81 == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_897); // @[FFT.scala 52:18]
  wire [31:0] _GEN_899 = 8'h82 == cnt[7:0] ? $signed(-32'shffec) : $signed(_GEN_898); // @[FFT.scala 52:18]
  wire [31:0] _GEN_900 = 8'h83 == cnt[7:0] ? $signed(-32'shffd4) : $signed(_GEN_899); // @[FFT.scala 52:18]
  wire [31:0] _GEN_901 = 8'h84 == cnt[7:0] ? $signed(-32'shffb1) : $signed(_GEN_900); // @[FFT.scala 52:18]
  wire [31:0] _GEN_902 = 8'h85 == cnt[7:0] ? $signed(-32'shff85) : $signed(_GEN_901); // @[FFT.scala 52:18]
  wire [31:0] _GEN_903 = 8'h86 == cnt[7:0] ? $signed(-32'shff4e) : $signed(_GEN_902); // @[FFT.scala 52:18]
  wire [31:0] _GEN_904 = 8'h87 == cnt[7:0] ? $signed(-32'shff0e) : $signed(_GEN_903); // @[FFT.scala 52:18]
  wire [31:0] _GEN_905 = 8'h88 == cnt[7:0] ? $signed(-32'shfec4) : $signed(_GEN_904); // @[FFT.scala 52:18]
  wire [31:0] _GEN_906 = 8'h89 == cnt[7:0] ? $signed(-32'shfe71) : $signed(_GEN_905); // @[FFT.scala 52:18]
  wire [31:0] _GEN_907 = 8'h8a == cnt[7:0] ? $signed(-32'shfe13) : $signed(_GEN_906); // @[FFT.scala 52:18]
  wire [31:0] _GEN_908 = 8'h8b == cnt[7:0] ? $signed(-32'shfdac) : $signed(_GEN_907); // @[FFT.scala 52:18]
  wire [31:0] _GEN_909 = 8'h8c == cnt[7:0] ? $signed(-32'shfd3b) : $signed(_GEN_908); // @[FFT.scala 52:18]
  wire [31:0] _GEN_910 = 8'h8d == cnt[7:0] ? $signed(-32'shfcc0) : $signed(_GEN_909); // @[FFT.scala 52:18]
  wire [31:0] _GEN_911 = 8'h8e == cnt[7:0] ? $signed(-32'shfc3b) : $signed(_GEN_910); // @[FFT.scala 52:18]
  wire [31:0] _GEN_912 = 8'h8f == cnt[7:0] ? $signed(-32'shfbad) : $signed(_GEN_911); // @[FFT.scala 52:18]
  wire [31:0] _GEN_913 = 8'h90 == cnt[7:0] ? $signed(-32'shfb15) : $signed(_GEN_912); // @[FFT.scala 52:18]
  wire [31:0] _GEN_914 = 8'h91 == cnt[7:0] ? $signed(-32'shfa73) : $signed(_GEN_913); // @[FFT.scala 52:18]
  wire [31:0] _GEN_915 = 8'h92 == cnt[7:0] ? $signed(-32'shf9c8) : $signed(_GEN_914); // @[FFT.scala 52:18]
  wire [31:0] _GEN_916 = 8'h93 == cnt[7:0] ? $signed(-32'shf913) : $signed(_GEN_915); // @[FFT.scala 52:18]
  wire [31:0] _GEN_917 = 8'h94 == cnt[7:0] ? $signed(-32'shf854) : $signed(_GEN_916); // @[FFT.scala 52:18]
  wire [31:0] _GEN_918 = 8'h95 == cnt[7:0] ? $signed(-32'shf78c) : $signed(_GEN_917); // @[FFT.scala 52:18]
  wire [31:0] _GEN_919 = 8'h96 == cnt[7:0] ? $signed(-32'shf6ba) : $signed(_GEN_918); // @[FFT.scala 52:18]
  wire [31:0] _GEN_920 = 8'h97 == cnt[7:0] ? $signed(-32'shf5df) : $signed(_GEN_919); // @[FFT.scala 52:18]
  wire [31:0] _GEN_921 = 8'h98 == cnt[7:0] ? $signed(-32'shf4fa) : $signed(_GEN_920); // @[FFT.scala 52:18]
  wire [31:0] _GEN_922 = 8'h99 == cnt[7:0] ? $signed(-32'shf40c) : $signed(_GEN_921); // @[FFT.scala 52:18]
  wire [31:0] _GEN_923 = 8'h9a == cnt[7:0] ? $signed(-32'shf314) : $signed(_GEN_922); // @[FFT.scala 52:18]
  wire [31:0] _GEN_924 = 8'h9b == cnt[7:0] ? $signed(-32'shf213) : $signed(_GEN_923); // @[FFT.scala 52:18]
  wire [31:0] _GEN_925 = 8'h9c == cnt[7:0] ? $signed(-32'shf109) : $signed(_GEN_924); // @[FFT.scala 52:18]
  wire [31:0] _GEN_926 = 8'h9d == cnt[7:0] ? $signed(-32'sheff5) : $signed(_GEN_925); // @[FFT.scala 52:18]
  wire [31:0] _GEN_927 = 8'h9e == cnt[7:0] ? $signed(-32'sheed9) : $signed(_GEN_926); // @[FFT.scala 52:18]
  wire [31:0] _GEN_928 = 8'h9f == cnt[7:0] ? $signed(-32'shedb3) : $signed(_GEN_927); // @[FFT.scala 52:18]
  wire [31:0] _GEN_929 = 8'ha0 == cnt[7:0] ? $signed(-32'shec83) : $signed(_GEN_928); // @[FFT.scala 52:18]
  wire [31:0] _GEN_930 = 8'ha1 == cnt[7:0] ? $signed(-32'sheb4b) : $signed(_GEN_929); // @[FFT.scala 52:18]
  wire [31:0] _GEN_931 = 8'ha2 == cnt[7:0] ? $signed(-32'shea0a) : $signed(_GEN_930); // @[FFT.scala 52:18]
  wire [31:0] _GEN_932 = 8'ha3 == cnt[7:0] ? $signed(-32'she8bf) : $signed(_GEN_931); // @[FFT.scala 52:18]
  wire [31:0] _GEN_933 = 8'ha4 == cnt[7:0] ? $signed(-32'she76c) : $signed(_GEN_932); // @[FFT.scala 52:18]
  wire [31:0] _GEN_934 = 8'ha5 == cnt[7:0] ? $signed(-32'she610) : $signed(_GEN_933); // @[FFT.scala 52:18]
  wire [31:0] _GEN_935 = 8'ha6 == cnt[7:0] ? $signed(-32'she4aa) : $signed(_GEN_934); // @[FFT.scala 52:18]
  wire [31:0] _GEN_936 = 8'ha7 == cnt[7:0] ? $signed(-32'she33c) : $signed(_GEN_935); // @[FFT.scala 52:18]
  wire [31:0] _GEN_937 = 8'ha8 == cnt[7:0] ? $signed(-32'she1c6) : $signed(_GEN_936); // @[FFT.scala 52:18]
  wire [31:0] _GEN_938 = 8'ha9 == cnt[7:0] ? $signed(-32'she046) : $signed(_GEN_937); // @[FFT.scala 52:18]
  wire [31:0] _GEN_939 = 8'haa == cnt[7:0] ? $signed(-32'shdebe) : $signed(_GEN_938); // @[FFT.scala 52:18]
  wire [31:0] _GEN_940 = 8'hab == cnt[7:0] ? $signed(-32'shdd2d) : $signed(_GEN_939); // @[FFT.scala 52:18]
  wire [31:0] _GEN_941 = 8'hac == cnt[7:0] ? $signed(-32'shdb94) : $signed(_GEN_940); // @[FFT.scala 52:18]
  wire [31:0] _GEN_942 = 8'had == cnt[7:0] ? $signed(-32'shd9f2) : $signed(_GEN_941); // @[FFT.scala 52:18]
  wire [31:0] _GEN_943 = 8'hae == cnt[7:0] ? $signed(-32'shd848) : $signed(_GEN_942); // @[FFT.scala 52:18]
  wire [31:0] _GEN_944 = 8'haf == cnt[7:0] ? $signed(-32'shd696) : $signed(_GEN_943); // @[FFT.scala 52:18]
  wire [31:0] _GEN_945 = 8'hb0 == cnt[7:0] ? $signed(-32'shd4db) : $signed(_GEN_944); // @[FFT.scala 52:18]
  wire [31:0] _GEN_946 = 8'hb1 == cnt[7:0] ? $signed(-32'shd318) : $signed(_GEN_945); // @[FFT.scala 52:18]
  wire [31:0] _GEN_947 = 8'hb2 == cnt[7:0] ? $signed(-32'shd14d) : $signed(_GEN_946); // @[FFT.scala 52:18]
  wire [31:0] _GEN_948 = 8'hb3 == cnt[7:0] ? $signed(-32'shcf7a) : $signed(_GEN_947); // @[FFT.scala 52:18]
  wire [31:0] _GEN_949 = 8'hb4 == cnt[7:0] ? $signed(-32'shcd9f) : $signed(_GEN_948); // @[FFT.scala 52:18]
  wire [31:0] _GEN_950 = 8'hb5 == cnt[7:0] ? $signed(-32'shcbbc) : $signed(_GEN_949); // @[FFT.scala 52:18]
  wire [31:0] _GEN_951 = 8'hb6 == cnt[7:0] ? $signed(-32'shc9d1) : $signed(_GEN_950); // @[FFT.scala 52:18]
  wire [31:0] _GEN_952 = 8'hb7 == cnt[7:0] ? $signed(-32'shc7de) : $signed(_GEN_951); // @[FFT.scala 52:18]
  wire [31:0] _GEN_953 = 8'hb8 == cnt[7:0] ? $signed(-32'shc5e4) : $signed(_GEN_952); // @[FFT.scala 52:18]
  wire [31:0] _GEN_954 = 8'hb9 == cnt[7:0] ? $signed(-32'shc3e2) : $signed(_GEN_953); // @[FFT.scala 52:18]
  wire [31:0] _GEN_955 = 8'hba == cnt[7:0] ? $signed(-32'shc1d8) : $signed(_GEN_954); // @[FFT.scala 52:18]
  wire [31:0] _GEN_956 = 8'hbb == cnt[7:0] ? $signed(-32'shbfc7) : $signed(_GEN_955); // @[FFT.scala 52:18]
  wire [31:0] _GEN_957 = 8'hbc == cnt[7:0] ? $signed(-32'shbdaf) : $signed(_GEN_956); // @[FFT.scala 52:18]
  wire [31:0] _GEN_958 = 8'hbd == cnt[7:0] ? $signed(-32'shbb8f) : $signed(_GEN_957); // @[FFT.scala 52:18]
  wire [31:0] _GEN_959 = 8'hbe == cnt[7:0] ? $signed(-32'shb968) : $signed(_GEN_958); // @[FFT.scala 52:18]
  wire [31:0] _GEN_960 = 8'hbf == cnt[7:0] ? $signed(-32'shb73a) : $signed(_GEN_959); // @[FFT.scala 52:18]
  wire [31:0] _GEN_961 = 8'hc0 == cnt[7:0] ? $signed(-32'shb505) : $signed(_GEN_960); // @[FFT.scala 52:18]
  wire [31:0] _GEN_962 = 8'hc1 == cnt[7:0] ? $signed(-32'shb2c9) : $signed(_GEN_961); // @[FFT.scala 52:18]
  wire [31:0] _GEN_963 = 8'hc2 == cnt[7:0] ? $signed(-32'shb086) : $signed(_GEN_962); // @[FFT.scala 52:18]
  wire [31:0] _GEN_964 = 8'hc3 == cnt[7:0] ? $signed(-32'shae3c) : $signed(_GEN_963); // @[FFT.scala 52:18]
  wire [31:0] _GEN_965 = 8'hc4 == cnt[7:0] ? $signed(-32'shabeb) : $signed(_GEN_964); // @[FFT.scala 52:18]
  wire [31:0] _GEN_966 = 8'hc5 == cnt[7:0] ? $signed(-32'sha994) : $signed(_GEN_965); // @[FFT.scala 52:18]
  wire [31:0] _GEN_967 = 8'hc6 == cnt[7:0] ? $signed(-32'sha736) : $signed(_GEN_966); // @[FFT.scala 52:18]
  wire [31:0] _GEN_968 = 8'hc7 == cnt[7:0] ? $signed(-32'sha4d2) : $signed(_GEN_967); // @[FFT.scala 52:18]
  wire [31:0] _GEN_969 = 8'hc8 == cnt[7:0] ? $signed(-32'sha268) : $signed(_GEN_968); // @[FFT.scala 52:18]
  wire [31:0] _GEN_970 = 8'hc9 == cnt[7:0] ? $signed(-32'sh9ff7) : $signed(_GEN_969); // @[FFT.scala 52:18]
  wire [31:0] _GEN_971 = 8'hca == cnt[7:0] ? $signed(-32'sh9d80) : $signed(_GEN_970); // @[FFT.scala 52:18]
  wire [31:0] _GEN_972 = 8'hcb == cnt[7:0] ? $signed(-32'sh9b03) : $signed(_GEN_971); // @[FFT.scala 52:18]
  wire [31:0] _GEN_973 = 8'hcc == cnt[7:0] ? $signed(-32'sh9880) : $signed(_GEN_972); // @[FFT.scala 52:18]
  wire [31:0] _GEN_974 = 8'hcd == cnt[7:0] ? $signed(-32'sh95f7) : $signed(_GEN_973); // @[FFT.scala 52:18]
  wire [31:0] _GEN_975 = 8'hce == cnt[7:0] ? $signed(-32'sh9368) : $signed(_GEN_974); // @[FFT.scala 52:18]
  wire [31:0] _GEN_976 = 8'hcf == cnt[7:0] ? $signed(-32'sh90d4) : $signed(_GEN_975); // @[FFT.scala 52:18]
  wire [31:0] _GEN_977 = 8'hd0 == cnt[7:0] ? $signed(-32'sh8e3a) : $signed(_GEN_976); // @[FFT.scala 52:18]
  wire [31:0] _GEN_978 = 8'hd1 == cnt[7:0] ? $signed(-32'sh8b9a) : $signed(_GEN_977); // @[FFT.scala 52:18]
  wire [31:0] _GEN_979 = 8'hd2 == cnt[7:0] ? $signed(-32'sh88f6) : $signed(_GEN_978); // @[FFT.scala 52:18]
  wire [31:0] _GEN_980 = 8'hd3 == cnt[7:0] ? $signed(-32'sh864c) : $signed(_GEN_979); // @[FFT.scala 52:18]
  wire [31:0] _GEN_981 = 8'hd4 == cnt[7:0] ? $signed(-32'sh839c) : $signed(_GEN_980); // @[FFT.scala 52:18]
  wire [31:0] _GEN_982 = 8'hd5 == cnt[7:0] ? $signed(-32'sh80e8) : $signed(_GEN_981); // @[FFT.scala 52:18]
  wire [31:0] _GEN_983 = 8'hd6 == cnt[7:0] ? $signed(-32'sh7e2f) : $signed(_GEN_982); // @[FFT.scala 52:18]
  wire [31:0] _GEN_984 = 8'hd7 == cnt[7:0] ? $signed(-32'sh7b70) : $signed(_GEN_983); // @[FFT.scala 52:18]
  wire [31:0] _GEN_985 = 8'hd8 == cnt[7:0] ? $signed(-32'sh78ad) : $signed(_GEN_984); // @[FFT.scala 52:18]
  wire [31:0] _GEN_986 = 8'hd9 == cnt[7:0] ? $signed(-32'sh75e6) : $signed(_GEN_985); // @[FFT.scala 52:18]
  wire [31:0] _GEN_987 = 8'hda == cnt[7:0] ? $signed(-32'sh731a) : $signed(_GEN_986); // @[FFT.scala 52:18]
  wire [31:0] _GEN_988 = 8'hdb == cnt[7:0] ? $signed(-32'sh7049) : $signed(_GEN_987); // @[FFT.scala 52:18]
  wire [31:0] _GEN_989 = 8'hdc == cnt[7:0] ? $signed(-32'sh6d74) : $signed(_GEN_988); // @[FFT.scala 52:18]
  wire [31:0] _GEN_990 = 8'hdd == cnt[7:0] ? $signed(-32'sh6a9b) : $signed(_GEN_989); // @[FFT.scala 52:18]
  wire [31:0] _GEN_991 = 8'hde == cnt[7:0] ? $signed(-32'sh67be) : $signed(_GEN_990); // @[FFT.scala 52:18]
  wire [31:0] _GEN_992 = 8'hdf == cnt[7:0] ? $signed(-32'sh64dd) : $signed(_GEN_991); // @[FFT.scala 52:18]
  wire [31:0] _GEN_993 = 8'he0 == cnt[7:0] ? $signed(-32'sh61f8) : $signed(_GEN_992); // @[FFT.scala 52:18]
  wire [31:0] _GEN_994 = 8'he1 == cnt[7:0] ? $signed(-32'sh5f0f) : $signed(_GEN_993); // @[FFT.scala 52:18]
  wire [31:0] _GEN_995 = 8'he2 == cnt[7:0] ? $signed(-32'sh5c22) : $signed(_GEN_994); // @[FFT.scala 52:18]
  wire [31:0] _GEN_996 = 8'he3 == cnt[7:0] ? $signed(-32'sh5932) : $signed(_GEN_995); // @[FFT.scala 52:18]
  wire [31:0] _GEN_997 = 8'he4 == cnt[7:0] ? $signed(-32'sh563e) : $signed(_GEN_996); // @[FFT.scala 52:18]
  wire [31:0] _GEN_998 = 8'he5 == cnt[7:0] ? $signed(-32'sh5348) : $signed(_GEN_997); // @[FFT.scala 52:18]
  wire [31:0] _GEN_999 = 8'he6 == cnt[7:0] ? $signed(-32'sh504d) : $signed(_GEN_998); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1000 = 8'he7 == cnt[7:0] ? $signed(-32'sh4d50) : $signed(_GEN_999); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1001 = 8'he8 == cnt[7:0] ? $signed(-32'sh4a50) : $signed(_GEN_1000); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1002 = 8'he9 == cnt[7:0] ? $signed(-32'sh474d) : $signed(_GEN_1001); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1003 = 8'hea == cnt[7:0] ? $signed(-32'sh4447) : $signed(_GEN_1002); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1004 = 8'heb == cnt[7:0] ? $signed(-32'sh413f) : $signed(_GEN_1003); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1005 = 8'hec == cnt[7:0] ? $signed(-32'sh3e34) : $signed(_GEN_1004); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1006 = 8'hed == cnt[7:0] ? $signed(-32'sh3b27) : $signed(_GEN_1005); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1007 = 8'hee == cnt[7:0] ? $signed(-32'sh3817) : $signed(_GEN_1006); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1008 = 8'hef == cnt[7:0] ? $signed(-32'sh3505) : $signed(_GEN_1007); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1009 = 8'hf0 == cnt[7:0] ? $signed(-32'sh31f1) : $signed(_GEN_1008); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1010 = 8'hf1 == cnt[7:0] ? $signed(-32'sh2edc) : $signed(_GEN_1009); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1011 = 8'hf2 == cnt[7:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1010); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1012 = 8'hf3 == cnt[7:0] ? $signed(-32'sh28ab) : $signed(_GEN_1011); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1013 = 8'hf4 == cnt[7:0] ? $signed(-32'sh2590) : $signed(_GEN_1012); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1014 = 8'hf5 == cnt[7:0] ? $signed(-32'sh2274) : $signed(_GEN_1013); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1015 = 8'hf6 == cnt[7:0] ? $signed(-32'sh1f56) : $signed(_GEN_1014); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1016 = 8'hf7 == cnt[7:0] ? $signed(-32'sh1c38) : $signed(_GEN_1015); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1017 = 8'hf8 == cnt[7:0] ? $signed(-32'sh1918) : $signed(_GEN_1016); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1018 = 8'hf9 == cnt[7:0] ? $signed(-32'sh15f7) : $signed(_GEN_1017); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1019 = 8'hfa == cnt[7:0] ? $signed(-32'sh12d5) : $signed(_GEN_1018); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1020 = 8'hfb == cnt[7:0] ? $signed(-32'shfb3) : $signed(_GEN_1019); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1021 = 8'hfc == cnt[7:0] ? $signed(-32'shc90) : $signed(_GEN_1020); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1022 = 8'hfd == cnt[7:0] ? $signed(-32'sh96c) : $signed(_GEN_1021); // @[FFT.scala 52:18]
  wire [31:0] _GEN_1023 = 8'hfe == cnt[7:0] ? $signed(-32'sh648) : $signed(_GEN_1022); // @[FFT.scala 52:18]
  reg [31:0] _T_150_re; // @[Reg.scala 15:16]
  reg [31:0] _T_150_im; // @[Reg.scala 15:16]
  reg [31:0] _T_151_re; // @[Reg.scala 15:16]
  reg [31:0] _T_151_im; // @[Reg.scala 15:16]
  reg [31:0] _T_152_re; // @[Reg.scala 15:16]
  reg [31:0] _T_152_im; // @[Reg.scala 15:16]
  reg [31:0] _T_153_re; // @[Reg.scala 15:16]
  reg [31:0] _T_153_im; // @[Reg.scala 15:16]
  reg [31:0] _T_154_re; // @[Reg.scala 15:16]
  reg [31:0] _T_154_im; // @[Reg.scala 15:16]
  reg [31:0] _T_155_re; // @[Reg.scala 15:16]
  reg [31:0] _T_155_im; // @[Reg.scala 15:16]
  reg [31:0] _T_156_re; // @[Reg.scala 15:16]
  reg [31:0] _T_156_im; // @[Reg.scala 15:16]
  reg [31:0] _T_157_re; // @[Reg.scala 15:16]
  reg [31:0] _T_157_im; // @[Reg.scala 15:16]
  reg [31:0] _T_158_re; // @[Reg.scala 15:16]
  reg [31:0] _T_158_im; // @[Reg.scala 15:16]
  reg [31:0] _T_159_re; // @[Reg.scala 15:16]
  reg [31:0] _T_159_im; // @[Reg.scala 15:16]
  reg [31:0] _T_160_re; // @[Reg.scala 15:16]
  reg [31:0] _T_160_im; // @[Reg.scala 15:16]
  reg [31:0] _T_161_re; // @[Reg.scala 15:16]
  reg [31:0] _T_161_im; // @[Reg.scala 15:16]
  reg [31:0] _T_162_re; // @[Reg.scala 15:16]
  reg [31:0] _T_162_im; // @[Reg.scala 15:16]
  reg [31:0] _T_163_re; // @[Reg.scala 15:16]
  reg [31:0] _T_163_im; // @[Reg.scala 15:16]
  reg [31:0] _T_164_re; // @[Reg.scala 15:16]
  reg [31:0] _T_164_im; // @[Reg.scala 15:16]
  reg [31:0] _T_165_re; // @[Reg.scala 15:16]
  reg [31:0] _T_165_im; // @[Reg.scala 15:16]
  reg [31:0] _T_166_re; // @[Reg.scala 15:16]
  reg [31:0] _T_166_im; // @[Reg.scala 15:16]
  reg [31:0] _T_167_re; // @[Reg.scala 15:16]
  reg [31:0] _T_167_im; // @[Reg.scala 15:16]
  reg [31:0] _T_168_re; // @[Reg.scala 15:16]
  reg [31:0] _T_168_im; // @[Reg.scala 15:16]
  reg [31:0] _T_169_re; // @[Reg.scala 15:16]
  reg [31:0] _T_169_im; // @[Reg.scala 15:16]
  reg [31:0] _T_170_re; // @[Reg.scala 15:16]
  reg [31:0] _T_170_im; // @[Reg.scala 15:16]
  reg [31:0] _T_171_re; // @[Reg.scala 15:16]
  reg [31:0] _T_171_im; // @[Reg.scala 15:16]
  reg [31:0] _T_172_re; // @[Reg.scala 15:16]
  reg [31:0] _T_172_im; // @[Reg.scala 15:16]
  reg [31:0] _T_173_re; // @[Reg.scala 15:16]
  reg [31:0] _T_173_im; // @[Reg.scala 15:16]
  reg [31:0] _T_174_re; // @[Reg.scala 15:16]
  reg [31:0] _T_174_im; // @[Reg.scala 15:16]
  reg [31:0] _T_175_re; // @[Reg.scala 15:16]
  reg [31:0] _T_175_im; // @[Reg.scala 15:16]
  reg [31:0] _T_176_re; // @[Reg.scala 15:16]
  reg [31:0] _T_176_im; // @[Reg.scala 15:16]
  reg [31:0] _T_177_re; // @[Reg.scala 15:16]
  reg [31:0] _T_177_im; // @[Reg.scala 15:16]
  reg [31:0] _T_178_re; // @[Reg.scala 15:16]
  reg [31:0] _T_178_im; // @[Reg.scala 15:16]
  reg [31:0] _T_179_re; // @[Reg.scala 15:16]
  reg [31:0] _T_179_im; // @[Reg.scala 15:16]
  reg [31:0] _T_180_re; // @[Reg.scala 15:16]
  reg [31:0] _T_180_im; // @[Reg.scala 15:16]
  reg [31:0] _T_181_re; // @[Reg.scala 15:16]
  reg [31:0] _T_181_im; // @[Reg.scala 15:16]
  reg [31:0] _T_182_re; // @[Reg.scala 15:16]
  reg [31:0] _T_182_im; // @[Reg.scala 15:16]
  reg [31:0] _T_183_re; // @[Reg.scala 15:16]
  reg [31:0] _T_183_im; // @[Reg.scala 15:16]
  reg [31:0] _T_184_re; // @[Reg.scala 15:16]
  reg [31:0] _T_184_im; // @[Reg.scala 15:16]
  reg [31:0] _T_185_re; // @[Reg.scala 15:16]
  reg [31:0] _T_185_im; // @[Reg.scala 15:16]
  reg [31:0] _T_186_re; // @[Reg.scala 15:16]
  reg [31:0] _T_186_im; // @[Reg.scala 15:16]
  reg [31:0] _T_187_re; // @[Reg.scala 15:16]
  reg [31:0] _T_187_im; // @[Reg.scala 15:16]
  reg [31:0] _T_188_re; // @[Reg.scala 15:16]
  reg [31:0] _T_188_im; // @[Reg.scala 15:16]
  reg [31:0] _T_189_re; // @[Reg.scala 15:16]
  reg [31:0] _T_189_im; // @[Reg.scala 15:16]
  reg [31:0] _T_190_re; // @[Reg.scala 15:16]
  reg [31:0] _T_190_im; // @[Reg.scala 15:16]
  reg [31:0] _T_191_re; // @[Reg.scala 15:16]
  reg [31:0] _T_191_im; // @[Reg.scala 15:16]
  reg [31:0] _T_192_re; // @[Reg.scala 15:16]
  reg [31:0] _T_192_im; // @[Reg.scala 15:16]
  reg [31:0] _T_193_re; // @[Reg.scala 15:16]
  reg [31:0] _T_193_im; // @[Reg.scala 15:16]
  reg [31:0] _T_194_re; // @[Reg.scala 15:16]
  reg [31:0] _T_194_im; // @[Reg.scala 15:16]
  reg [31:0] _T_195_re; // @[Reg.scala 15:16]
  reg [31:0] _T_195_im; // @[Reg.scala 15:16]
  reg [31:0] _T_196_re; // @[Reg.scala 15:16]
  reg [31:0] _T_196_im; // @[Reg.scala 15:16]
  reg [31:0] _T_197_re; // @[Reg.scala 15:16]
  reg [31:0] _T_197_im; // @[Reg.scala 15:16]
  reg [31:0] _T_198_re; // @[Reg.scala 15:16]
  reg [31:0] _T_198_im; // @[Reg.scala 15:16]
  reg [31:0] _T_199_re; // @[Reg.scala 15:16]
  reg [31:0] _T_199_im; // @[Reg.scala 15:16]
  reg [31:0] _T_200_re; // @[Reg.scala 15:16]
  reg [31:0] _T_200_im; // @[Reg.scala 15:16]
  reg [31:0] _T_201_re; // @[Reg.scala 15:16]
  reg [31:0] _T_201_im; // @[Reg.scala 15:16]
  reg [31:0] _T_202_re; // @[Reg.scala 15:16]
  reg [31:0] _T_202_im; // @[Reg.scala 15:16]
  reg [31:0] _T_203_re; // @[Reg.scala 15:16]
  reg [31:0] _T_203_im; // @[Reg.scala 15:16]
  reg [31:0] _T_204_re; // @[Reg.scala 15:16]
  reg [31:0] _T_204_im; // @[Reg.scala 15:16]
  reg [31:0] _T_205_re; // @[Reg.scala 15:16]
  reg [31:0] _T_205_im; // @[Reg.scala 15:16]
  reg [31:0] _T_206_re; // @[Reg.scala 15:16]
  reg [31:0] _T_206_im; // @[Reg.scala 15:16]
  reg [31:0] _T_207_re; // @[Reg.scala 15:16]
  reg [31:0] _T_207_im; // @[Reg.scala 15:16]
  reg [31:0] _T_208_re; // @[Reg.scala 15:16]
  reg [31:0] _T_208_im; // @[Reg.scala 15:16]
  reg [31:0] _T_209_re; // @[Reg.scala 15:16]
  reg [31:0] _T_209_im; // @[Reg.scala 15:16]
  reg [31:0] _T_210_re; // @[Reg.scala 15:16]
  reg [31:0] _T_210_im; // @[Reg.scala 15:16]
  reg [31:0] _T_211_re; // @[Reg.scala 15:16]
  reg [31:0] _T_211_im; // @[Reg.scala 15:16]
  reg [31:0] _T_212_re; // @[Reg.scala 15:16]
  reg [31:0] _T_212_im; // @[Reg.scala 15:16]
  reg [31:0] _T_213_re; // @[Reg.scala 15:16]
  reg [31:0] _T_213_im; // @[Reg.scala 15:16]
  reg [31:0] _T_214_re; // @[Reg.scala 15:16]
  reg [31:0] _T_214_im; // @[Reg.scala 15:16]
  reg [31:0] _T_215_re; // @[Reg.scala 15:16]
  reg [31:0] _T_215_im; // @[Reg.scala 15:16]
  reg [31:0] _T_216_re; // @[Reg.scala 15:16]
  reg [31:0] _T_216_im; // @[Reg.scala 15:16]
  reg [31:0] _T_217_re; // @[Reg.scala 15:16]
  reg [31:0] _T_217_im; // @[Reg.scala 15:16]
  reg [31:0] _T_218_re; // @[Reg.scala 15:16]
  reg [31:0] _T_218_im; // @[Reg.scala 15:16]
  reg [31:0] _T_219_re; // @[Reg.scala 15:16]
  reg [31:0] _T_219_im; // @[Reg.scala 15:16]
  reg [31:0] _T_220_re; // @[Reg.scala 15:16]
  reg [31:0] _T_220_im; // @[Reg.scala 15:16]
  reg [31:0] _T_221_re; // @[Reg.scala 15:16]
  reg [31:0] _T_221_im; // @[Reg.scala 15:16]
  reg [31:0] _T_222_re; // @[Reg.scala 15:16]
  reg [31:0] _T_222_im; // @[Reg.scala 15:16]
  reg [31:0] _T_223_re; // @[Reg.scala 15:16]
  reg [31:0] _T_223_im; // @[Reg.scala 15:16]
  reg [31:0] _T_224_re; // @[Reg.scala 15:16]
  reg [31:0] _T_224_im; // @[Reg.scala 15:16]
  reg [31:0] _T_225_re; // @[Reg.scala 15:16]
  reg [31:0] _T_225_im; // @[Reg.scala 15:16]
  reg [31:0] _T_226_re; // @[Reg.scala 15:16]
  reg [31:0] _T_226_im; // @[Reg.scala 15:16]
  reg [31:0] _T_227_re; // @[Reg.scala 15:16]
  reg [31:0] _T_227_im; // @[Reg.scala 15:16]
  reg [31:0] _T_228_re; // @[Reg.scala 15:16]
  reg [31:0] _T_228_im; // @[Reg.scala 15:16]
  reg [31:0] _T_229_re; // @[Reg.scala 15:16]
  reg [31:0] _T_229_im; // @[Reg.scala 15:16]
  reg [31:0] _T_230_re; // @[Reg.scala 15:16]
  reg [31:0] _T_230_im; // @[Reg.scala 15:16]
  reg [31:0] _T_231_re; // @[Reg.scala 15:16]
  reg [31:0] _T_231_im; // @[Reg.scala 15:16]
  reg [31:0] _T_232_re; // @[Reg.scala 15:16]
  reg [31:0] _T_232_im; // @[Reg.scala 15:16]
  reg [31:0] _T_233_re; // @[Reg.scala 15:16]
  reg [31:0] _T_233_im; // @[Reg.scala 15:16]
  reg [31:0] _T_234_re; // @[Reg.scala 15:16]
  reg [31:0] _T_234_im; // @[Reg.scala 15:16]
  reg [31:0] _T_235_re; // @[Reg.scala 15:16]
  reg [31:0] _T_235_im; // @[Reg.scala 15:16]
  reg [31:0] _T_236_re; // @[Reg.scala 15:16]
  reg [31:0] _T_236_im; // @[Reg.scala 15:16]
  reg [31:0] _T_237_re; // @[Reg.scala 15:16]
  reg [31:0] _T_237_im; // @[Reg.scala 15:16]
  reg [31:0] _T_238_re; // @[Reg.scala 15:16]
  reg [31:0] _T_238_im; // @[Reg.scala 15:16]
  reg [31:0] _T_239_re; // @[Reg.scala 15:16]
  reg [31:0] _T_239_im; // @[Reg.scala 15:16]
  reg [31:0] _T_240_re; // @[Reg.scala 15:16]
  reg [31:0] _T_240_im; // @[Reg.scala 15:16]
  reg [31:0] _T_241_re; // @[Reg.scala 15:16]
  reg [31:0] _T_241_im; // @[Reg.scala 15:16]
  reg [31:0] _T_242_re; // @[Reg.scala 15:16]
  reg [31:0] _T_242_im; // @[Reg.scala 15:16]
  reg [31:0] _T_243_re; // @[Reg.scala 15:16]
  reg [31:0] _T_243_im; // @[Reg.scala 15:16]
  reg [31:0] _T_244_re; // @[Reg.scala 15:16]
  reg [31:0] _T_244_im; // @[Reg.scala 15:16]
  reg [31:0] _T_245_re; // @[Reg.scala 15:16]
  reg [31:0] _T_245_im; // @[Reg.scala 15:16]
  reg [31:0] _T_246_re; // @[Reg.scala 15:16]
  reg [31:0] _T_246_im; // @[Reg.scala 15:16]
  reg [31:0] _T_247_re; // @[Reg.scala 15:16]
  reg [31:0] _T_247_im; // @[Reg.scala 15:16]
  reg [31:0] _T_248_re; // @[Reg.scala 15:16]
  reg [31:0] _T_248_im; // @[Reg.scala 15:16]
  reg [31:0] _T_249_re; // @[Reg.scala 15:16]
  reg [31:0] _T_249_im; // @[Reg.scala 15:16]
  reg [31:0] _T_250_re; // @[Reg.scala 15:16]
  reg [31:0] _T_250_im; // @[Reg.scala 15:16]
  reg [31:0] _T_251_re; // @[Reg.scala 15:16]
  reg [31:0] _T_251_im; // @[Reg.scala 15:16]
  reg [31:0] _T_252_re; // @[Reg.scala 15:16]
  reg [31:0] _T_252_im; // @[Reg.scala 15:16]
  reg [31:0] _T_253_re; // @[Reg.scala 15:16]
  reg [31:0] _T_253_im; // @[Reg.scala 15:16]
  reg [31:0] _T_254_re; // @[Reg.scala 15:16]
  reg [31:0] _T_254_im; // @[Reg.scala 15:16]
  reg [31:0] _T_255_re; // @[Reg.scala 15:16]
  reg [31:0] _T_255_im; // @[Reg.scala 15:16]
  reg [31:0] _T_256_re; // @[Reg.scala 15:16]
  reg [31:0] _T_256_im; // @[Reg.scala 15:16]
  reg [31:0] _T_257_re; // @[Reg.scala 15:16]
  reg [31:0] _T_257_im; // @[Reg.scala 15:16]
  reg [31:0] _T_258_re; // @[Reg.scala 15:16]
  reg [31:0] _T_258_im; // @[Reg.scala 15:16]
  reg [31:0] _T_259_re; // @[Reg.scala 15:16]
  reg [31:0] _T_259_im; // @[Reg.scala 15:16]
  reg [31:0] _T_260_re; // @[Reg.scala 15:16]
  reg [31:0] _T_260_im; // @[Reg.scala 15:16]
  reg [31:0] _T_261_re; // @[Reg.scala 15:16]
  reg [31:0] _T_261_im; // @[Reg.scala 15:16]
  reg [31:0] _T_262_re; // @[Reg.scala 15:16]
  reg [31:0] _T_262_im; // @[Reg.scala 15:16]
  reg [31:0] _T_263_re; // @[Reg.scala 15:16]
  reg [31:0] _T_263_im; // @[Reg.scala 15:16]
  reg [31:0] _T_264_re; // @[Reg.scala 15:16]
  reg [31:0] _T_264_im; // @[Reg.scala 15:16]
  reg [31:0] _T_265_re; // @[Reg.scala 15:16]
  reg [31:0] _T_265_im; // @[Reg.scala 15:16]
  reg [31:0] _T_266_re; // @[Reg.scala 15:16]
  reg [31:0] _T_266_im; // @[Reg.scala 15:16]
  reg [31:0] _T_267_re; // @[Reg.scala 15:16]
  reg [31:0] _T_267_im; // @[Reg.scala 15:16]
  reg [31:0] _T_268_re; // @[Reg.scala 15:16]
  reg [31:0] _T_268_im; // @[Reg.scala 15:16]
  reg [31:0] _T_269_re; // @[Reg.scala 15:16]
  reg [31:0] _T_269_im; // @[Reg.scala 15:16]
  reg [31:0] _T_270_re; // @[Reg.scala 15:16]
  reg [31:0] _T_270_im; // @[Reg.scala 15:16]
  reg [31:0] _T_271_re; // @[Reg.scala 15:16]
  reg [31:0] _T_271_im; // @[Reg.scala 15:16]
  reg [31:0] _T_272_re; // @[Reg.scala 15:16]
  reg [31:0] _T_272_im; // @[Reg.scala 15:16]
  reg [31:0] _T_273_re; // @[Reg.scala 15:16]
  reg [31:0] _T_273_im; // @[Reg.scala 15:16]
  reg [31:0] _T_274_re; // @[Reg.scala 15:16]
  reg [31:0] _T_274_im; // @[Reg.scala 15:16]
  reg [31:0] _T_275_re; // @[Reg.scala 15:16]
  reg [31:0] _T_275_im; // @[Reg.scala 15:16]
  reg [31:0] _T_276_re; // @[Reg.scala 15:16]
  reg [31:0] _T_276_im; // @[Reg.scala 15:16]
  reg [31:0] _T_277_re; // @[Reg.scala 15:16]
  reg [31:0] _T_277_im; // @[Reg.scala 15:16]
  reg [31:0] _T_278_re; // @[Reg.scala 15:16]
  reg [31:0] _T_278_im; // @[Reg.scala 15:16]
  reg [31:0] _T_279_re; // @[Reg.scala 15:16]
  reg [31:0] _T_279_im; // @[Reg.scala 15:16]
  reg [31:0] _T_280_re; // @[Reg.scala 15:16]
  reg [31:0] _T_280_im; // @[Reg.scala 15:16]
  reg [31:0] _T_281_re; // @[Reg.scala 15:16]
  reg [31:0] _T_281_im; // @[Reg.scala 15:16]
  reg [31:0] _T_282_re; // @[Reg.scala 15:16]
  reg [31:0] _T_282_im; // @[Reg.scala 15:16]
  reg [31:0] _T_283_re; // @[Reg.scala 15:16]
  reg [31:0] _T_283_im; // @[Reg.scala 15:16]
  reg [31:0] _T_284_re; // @[Reg.scala 15:16]
  reg [31:0] _T_284_im; // @[Reg.scala 15:16]
  reg [31:0] _T_285_re; // @[Reg.scala 15:16]
  reg [31:0] _T_285_im; // @[Reg.scala 15:16]
  reg [31:0] _T_286_re; // @[Reg.scala 15:16]
  reg [31:0] _T_286_im; // @[Reg.scala 15:16]
  reg [31:0] _T_287_re; // @[Reg.scala 15:16]
  reg [31:0] _T_287_im; // @[Reg.scala 15:16]
  reg [31:0] _T_288_re; // @[Reg.scala 15:16]
  reg [31:0] _T_288_im; // @[Reg.scala 15:16]
  reg [31:0] _T_289_re; // @[Reg.scala 15:16]
  reg [31:0] _T_289_im; // @[Reg.scala 15:16]
  reg [31:0] _T_290_re; // @[Reg.scala 15:16]
  reg [31:0] _T_290_im; // @[Reg.scala 15:16]
  reg [31:0] _T_291_re; // @[Reg.scala 15:16]
  reg [31:0] _T_291_im; // @[Reg.scala 15:16]
  reg [31:0] _T_292_re; // @[Reg.scala 15:16]
  reg [31:0] _T_292_im; // @[Reg.scala 15:16]
  reg [31:0] _T_293_re; // @[Reg.scala 15:16]
  reg [31:0] _T_293_im; // @[Reg.scala 15:16]
  reg [31:0] _T_294_re; // @[Reg.scala 15:16]
  reg [31:0] _T_294_im; // @[Reg.scala 15:16]
  reg [31:0] _T_295_re; // @[Reg.scala 15:16]
  reg [31:0] _T_295_im; // @[Reg.scala 15:16]
  reg [31:0] _T_296_re; // @[Reg.scala 15:16]
  reg [31:0] _T_296_im; // @[Reg.scala 15:16]
  reg [31:0] _T_297_re; // @[Reg.scala 15:16]
  reg [31:0] _T_297_im; // @[Reg.scala 15:16]
  reg [31:0] _T_298_re; // @[Reg.scala 15:16]
  reg [31:0] _T_298_im; // @[Reg.scala 15:16]
  reg [31:0] _T_299_re; // @[Reg.scala 15:16]
  reg [31:0] _T_299_im; // @[Reg.scala 15:16]
  reg [31:0] _T_300_re; // @[Reg.scala 15:16]
  reg [31:0] _T_300_im; // @[Reg.scala 15:16]
  reg [31:0] _T_301_re; // @[Reg.scala 15:16]
  reg [31:0] _T_301_im; // @[Reg.scala 15:16]
  reg [31:0] _T_302_re; // @[Reg.scala 15:16]
  reg [31:0] _T_302_im; // @[Reg.scala 15:16]
  reg [31:0] _T_303_re; // @[Reg.scala 15:16]
  reg [31:0] _T_303_im; // @[Reg.scala 15:16]
  reg [31:0] _T_304_re; // @[Reg.scala 15:16]
  reg [31:0] _T_304_im; // @[Reg.scala 15:16]
  reg [31:0] _T_305_re; // @[Reg.scala 15:16]
  reg [31:0] _T_305_im; // @[Reg.scala 15:16]
  reg [31:0] _T_306_re; // @[Reg.scala 15:16]
  reg [31:0] _T_306_im; // @[Reg.scala 15:16]
  reg [31:0] _T_307_re; // @[Reg.scala 15:16]
  reg [31:0] _T_307_im; // @[Reg.scala 15:16]
  reg [31:0] _T_308_re; // @[Reg.scala 15:16]
  reg [31:0] _T_308_im; // @[Reg.scala 15:16]
  reg [31:0] _T_309_re; // @[Reg.scala 15:16]
  reg [31:0] _T_309_im; // @[Reg.scala 15:16]
  reg [31:0] _T_310_re; // @[Reg.scala 15:16]
  reg [31:0] _T_310_im; // @[Reg.scala 15:16]
  reg [31:0] _T_311_re; // @[Reg.scala 15:16]
  reg [31:0] _T_311_im; // @[Reg.scala 15:16]
  reg [31:0] _T_312_re; // @[Reg.scala 15:16]
  reg [31:0] _T_312_im; // @[Reg.scala 15:16]
  reg [31:0] _T_313_re; // @[Reg.scala 15:16]
  reg [31:0] _T_313_im; // @[Reg.scala 15:16]
  reg [31:0] _T_314_re; // @[Reg.scala 15:16]
  reg [31:0] _T_314_im; // @[Reg.scala 15:16]
  reg [31:0] _T_315_re; // @[Reg.scala 15:16]
  reg [31:0] _T_315_im; // @[Reg.scala 15:16]
  reg [31:0] _T_316_re; // @[Reg.scala 15:16]
  reg [31:0] _T_316_im; // @[Reg.scala 15:16]
  reg [31:0] _T_317_re; // @[Reg.scala 15:16]
  reg [31:0] _T_317_im; // @[Reg.scala 15:16]
  reg [31:0] _T_318_re; // @[Reg.scala 15:16]
  reg [31:0] _T_318_im; // @[Reg.scala 15:16]
  reg [31:0] _T_319_re; // @[Reg.scala 15:16]
  reg [31:0] _T_319_im; // @[Reg.scala 15:16]
  reg [31:0] _T_320_re; // @[Reg.scala 15:16]
  reg [31:0] _T_320_im; // @[Reg.scala 15:16]
  reg [31:0] _T_321_re; // @[Reg.scala 15:16]
  reg [31:0] _T_321_im; // @[Reg.scala 15:16]
  reg [31:0] _T_322_re; // @[Reg.scala 15:16]
  reg [31:0] _T_322_im; // @[Reg.scala 15:16]
  reg [31:0] _T_323_re; // @[Reg.scala 15:16]
  reg [31:0] _T_323_im; // @[Reg.scala 15:16]
  reg [31:0] _T_324_re; // @[Reg.scala 15:16]
  reg [31:0] _T_324_im; // @[Reg.scala 15:16]
  reg [31:0] _T_325_re; // @[Reg.scala 15:16]
  reg [31:0] _T_325_im; // @[Reg.scala 15:16]
  reg [31:0] _T_326_re; // @[Reg.scala 15:16]
  reg [31:0] _T_326_im; // @[Reg.scala 15:16]
  reg [31:0] _T_327_re; // @[Reg.scala 15:16]
  reg [31:0] _T_327_im; // @[Reg.scala 15:16]
  reg [31:0] _T_328_re; // @[Reg.scala 15:16]
  reg [31:0] _T_328_im; // @[Reg.scala 15:16]
  reg [31:0] _T_329_re; // @[Reg.scala 15:16]
  reg [31:0] _T_329_im; // @[Reg.scala 15:16]
  reg [31:0] _T_330_re; // @[Reg.scala 15:16]
  reg [31:0] _T_330_im; // @[Reg.scala 15:16]
  reg [31:0] _T_331_re; // @[Reg.scala 15:16]
  reg [31:0] _T_331_im; // @[Reg.scala 15:16]
  reg [31:0] _T_332_re; // @[Reg.scala 15:16]
  reg [31:0] _T_332_im; // @[Reg.scala 15:16]
  reg [31:0] _T_333_re; // @[Reg.scala 15:16]
  reg [31:0] _T_333_im; // @[Reg.scala 15:16]
  reg [31:0] _T_334_re; // @[Reg.scala 15:16]
  reg [31:0] _T_334_im; // @[Reg.scala 15:16]
  reg [31:0] _T_335_re; // @[Reg.scala 15:16]
  reg [31:0] _T_335_im; // @[Reg.scala 15:16]
  reg [31:0] _T_336_re; // @[Reg.scala 15:16]
  reg [31:0] _T_336_im; // @[Reg.scala 15:16]
  reg [31:0] _T_337_re; // @[Reg.scala 15:16]
  reg [31:0] _T_337_im; // @[Reg.scala 15:16]
  reg [31:0] _T_338_re; // @[Reg.scala 15:16]
  reg [31:0] _T_338_im; // @[Reg.scala 15:16]
  reg [31:0] _T_339_re; // @[Reg.scala 15:16]
  reg [31:0] _T_339_im; // @[Reg.scala 15:16]
  reg [31:0] _T_340_re; // @[Reg.scala 15:16]
  reg [31:0] _T_340_im; // @[Reg.scala 15:16]
  reg [31:0] _T_341_re; // @[Reg.scala 15:16]
  reg [31:0] _T_341_im; // @[Reg.scala 15:16]
  reg [31:0] _T_342_re; // @[Reg.scala 15:16]
  reg [31:0] _T_342_im; // @[Reg.scala 15:16]
  reg [31:0] _T_343_re; // @[Reg.scala 15:16]
  reg [31:0] _T_343_im; // @[Reg.scala 15:16]
  reg [31:0] _T_344_re; // @[Reg.scala 15:16]
  reg [31:0] _T_344_im; // @[Reg.scala 15:16]
  reg [31:0] _T_345_re; // @[Reg.scala 15:16]
  reg [31:0] _T_345_im; // @[Reg.scala 15:16]
  reg [31:0] _T_346_re; // @[Reg.scala 15:16]
  reg [31:0] _T_346_im; // @[Reg.scala 15:16]
  reg [31:0] _T_347_re; // @[Reg.scala 15:16]
  reg [31:0] _T_347_im; // @[Reg.scala 15:16]
  reg [31:0] _T_348_re; // @[Reg.scala 15:16]
  reg [31:0] _T_348_im; // @[Reg.scala 15:16]
  reg [31:0] _T_349_re; // @[Reg.scala 15:16]
  reg [31:0] _T_349_im; // @[Reg.scala 15:16]
  reg [31:0] _T_350_re; // @[Reg.scala 15:16]
  reg [31:0] _T_350_im; // @[Reg.scala 15:16]
  reg [31:0] _T_351_re; // @[Reg.scala 15:16]
  reg [31:0] _T_351_im; // @[Reg.scala 15:16]
  reg [31:0] _T_352_re; // @[Reg.scala 15:16]
  reg [31:0] _T_352_im; // @[Reg.scala 15:16]
  reg [31:0] _T_353_re; // @[Reg.scala 15:16]
  reg [31:0] _T_353_im; // @[Reg.scala 15:16]
  reg [31:0] _T_354_re; // @[Reg.scala 15:16]
  reg [31:0] _T_354_im; // @[Reg.scala 15:16]
  reg [31:0] _T_355_re; // @[Reg.scala 15:16]
  reg [31:0] _T_355_im; // @[Reg.scala 15:16]
  reg [31:0] _T_356_re; // @[Reg.scala 15:16]
  reg [31:0] _T_356_im; // @[Reg.scala 15:16]
  reg [31:0] _T_357_re; // @[Reg.scala 15:16]
  reg [31:0] _T_357_im; // @[Reg.scala 15:16]
  reg [31:0] _T_358_re; // @[Reg.scala 15:16]
  reg [31:0] _T_358_im; // @[Reg.scala 15:16]
  reg [31:0] _T_359_re; // @[Reg.scala 15:16]
  reg [31:0] _T_359_im; // @[Reg.scala 15:16]
  reg [31:0] _T_360_re; // @[Reg.scala 15:16]
  reg [31:0] _T_360_im; // @[Reg.scala 15:16]
  reg [31:0] _T_361_re; // @[Reg.scala 15:16]
  reg [31:0] _T_361_im; // @[Reg.scala 15:16]
  reg [31:0] _T_362_re; // @[Reg.scala 15:16]
  reg [31:0] _T_362_im; // @[Reg.scala 15:16]
  reg [31:0] _T_363_re; // @[Reg.scala 15:16]
  reg [31:0] _T_363_im; // @[Reg.scala 15:16]
  reg [31:0] _T_364_re; // @[Reg.scala 15:16]
  reg [31:0] _T_364_im; // @[Reg.scala 15:16]
  reg [31:0] _T_365_re; // @[Reg.scala 15:16]
  reg [31:0] _T_365_im; // @[Reg.scala 15:16]
  reg [31:0] _T_366_re; // @[Reg.scala 15:16]
  reg [31:0] _T_366_im; // @[Reg.scala 15:16]
  reg [31:0] _T_367_re; // @[Reg.scala 15:16]
  reg [31:0] _T_367_im; // @[Reg.scala 15:16]
  reg [31:0] _T_368_re; // @[Reg.scala 15:16]
  reg [31:0] _T_368_im; // @[Reg.scala 15:16]
  reg [31:0] _T_369_re; // @[Reg.scala 15:16]
  reg [31:0] _T_369_im; // @[Reg.scala 15:16]
  reg [31:0] _T_370_re; // @[Reg.scala 15:16]
  reg [31:0] _T_370_im; // @[Reg.scala 15:16]
  reg [31:0] _T_371_re; // @[Reg.scala 15:16]
  reg [31:0] _T_371_im; // @[Reg.scala 15:16]
  reg [31:0] _T_372_re; // @[Reg.scala 15:16]
  reg [31:0] _T_372_im; // @[Reg.scala 15:16]
  reg [31:0] _T_373_re; // @[Reg.scala 15:16]
  reg [31:0] _T_373_im; // @[Reg.scala 15:16]
  reg [31:0] _T_374_re; // @[Reg.scala 15:16]
  reg [31:0] _T_374_im; // @[Reg.scala 15:16]
  reg [31:0] _T_375_re; // @[Reg.scala 15:16]
  reg [31:0] _T_375_im; // @[Reg.scala 15:16]
  reg [31:0] _T_376_re; // @[Reg.scala 15:16]
  reg [31:0] _T_376_im; // @[Reg.scala 15:16]
  reg [31:0] _T_377_re; // @[Reg.scala 15:16]
  reg [31:0] _T_377_im; // @[Reg.scala 15:16]
  reg [31:0] _T_378_re; // @[Reg.scala 15:16]
  reg [31:0] _T_378_im; // @[Reg.scala 15:16]
  reg [31:0] _T_379_re; // @[Reg.scala 15:16]
  reg [31:0] _T_379_im; // @[Reg.scala 15:16]
  reg [31:0] _T_380_re; // @[Reg.scala 15:16]
  reg [31:0] _T_380_im; // @[Reg.scala 15:16]
  reg [31:0] _T_381_re; // @[Reg.scala 15:16]
  reg [31:0] _T_381_im; // @[Reg.scala 15:16]
  reg [31:0] _T_382_re; // @[Reg.scala 15:16]
  reg [31:0] _T_382_im; // @[Reg.scala 15:16]
  reg [31:0] _T_383_re; // @[Reg.scala 15:16]
  reg [31:0] _T_383_im; // @[Reg.scala 15:16]
  reg [31:0] _T_384_re; // @[Reg.scala 15:16]
  reg [31:0] _T_384_im; // @[Reg.scala 15:16]
  reg [31:0] _T_385_re; // @[Reg.scala 15:16]
  reg [31:0] _T_385_im; // @[Reg.scala 15:16]
  reg [31:0] _T_386_re; // @[Reg.scala 15:16]
  reg [31:0] _T_386_im; // @[Reg.scala 15:16]
  reg [31:0] _T_387_re; // @[Reg.scala 15:16]
  reg [31:0] _T_387_im; // @[Reg.scala 15:16]
  reg [31:0] _T_388_re; // @[Reg.scala 15:16]
  reg [31:0] _T_388_im; // @[Reg.scala 15:16]
  reg [31:0] _T_389_re; // @[Reg.scala 15:16]
  reg [31:0] _T_389_im; // @[Reg.scala 15:16]
  reg [31:0] _T_390_re; // @[Reg.scala 15:16]
  reg [31:0] _T_390_im; // @[Reg.scala 15:16]
  reg [31:0] _T_391_re; // @[Reg.scala 15:16]
  reg [31:0] _T_391_im; // @[Reg.scala 15:16]
  reg [31:0] _T_392_re; // @[Reg.scala 15:16]
  reg [31:0] _T_392_im; // @[Reg.scala 15:16]
  reg [31:0] _T_393_re; // @[Reg.scala 15:16]
  reg [31:0] _T_393_im; // @[Reg.scala 15:16]
  reg [31:0] _T_394_re; // @[Reg.scala 15:16]
  reg [31:0] _T_394_im; // @[Reg.scala 15:16]
  reg [31:0] _T_395_re; // @[Reg.scala 15:16]
  reg [31:0] _T_395_im; // @[Reg.scala 15:16]
  reg [31:0] _T_396_re; // @[Reg.scala 15:16]
  reg [31:0] _T_396_im; // @[Reg.scala 15:16]
  reg [31:0] _T_397_re; // @[Reg.scala 15:16]
  reg [31:0] _T_397_im; // @[Reg.scala 15:16]
  reg [31:0] _T_398_re; // @[Reg.scala 15:16]
  reg [31:0] _T_398_im; // @[Reg.scala 15:16]
  reg [31:0] _T_399_re; // @[Reg.scala 15:16]
  reg [31:0] _T_399_im; // @[Reg.scala 15:16]
  reg [31:0] _T_400_re; // @[Reg.scala 15:16]
  reg [31:0] _T_400_im; // @[Reg.scala 15:16]
  reg [31:0] _T_401_re; // @[Reg.scala 15:16]
  reg [31:0] _T_401_im; // @[Reg.scala 15:16]
  reg [31:0] _T_402_re; // @[Reg.scala 15:16]
  reg [31:0] _T_402_im; // @[Reg.scala 15:16]
  reg [31:0] _T_403_re; // @[Reg.scala 15:16]
  reg [31:0] _T_403_im; // @[Reg.scala 15:16]
  reg [31:0] _T_404_re; // @[Reg.scala 15:16]
  reg [31:0] _T_404_im; // @[Reg.scala 15:16]
  reg [31:0] _T_405_re; // @[Reg.scala 15:16]
  reg [31:0] _T_405_im; // @[Reg.scala 15:16]
  reg [31:0] _T_407_re; // @[Reg.scala 15:16]
  reg [31:0] _T_407_im; // @[Reg.scala 15:16]
  reg [31:0] _T_408_re; // @[Reg.scala 15:16]
  reg [31:0] _T_408_im; // @[Reg.scala 15:16]
  reg [31:0] _T_409_re; // @[Reg.scala 15:16]
  reg [31:0] _T_409_im; // @[Reg.scala 15:16]
  reg [31:0] _T_410_re; // @[Reg.scala 15:16]
  reg [31:0] _T_410_im; // @[Reg.scala 15:16]
  reg [31:0] _T_411_re; // @[Reg.scala 15:16]
  reg [31:0] _T_411_im; // @[Reg.scala 15:16]
  reg [31:0] _T_412_re; // @[Reg.scala 15:16]
  reg [31:0] _T_412_im; // @[Reg.scala 15:16]
  reg [31:0] _T_413_re; // @[Reg.scala 15:16]
  reg [31:0] _T_413_im; // @[Reg.scala 15:16]
  reg [31:0] _T_414_re; // @[Reg.scala 15:16]
  reg [31:0] _T_414_im; // @[Reg.scala 15:16]
  reg [31:0] _T_415_re; // @[Reg.scala 15:16]
  reg [31:0] _T_415_im; // @[Reg.scala 15:16]
  reg [31:0] _T_416_re; // @[Reg.scala 15:16]
  reg [31:0] _T_416_im; // @[Reg.scala 15:16]
  reg [31:0] _T_417_re; // @[Reg.scala 15:16]
  reg [31:0] _T_417_im; // @[Reg.scala 15:16]
  reg [31:0] _T_418_re; // @[Reg.scala 15:16]
  reg [31:0] _T_418_im; // @[Reg.scala 15:16]
  reg [31:0] _T_419_re; // @[Reg.scala 15:16]
  reg [31:0] _T_419_im; // @[Reg.scala 15:16]
  reg [31:0] _T_420_re; // @[Reg.scala 15:16]
  reg [31:0] _T_420_im; // @[Reg.scala 15:16]
  reg [31:0] _T_421_re; // @[Reg.scala 15:16]
  reg [31:0] _T_421_im; // @[Reg.scala 15:16]
  reg [31:0] _T_422_re; // @[Reg.scala 15:16]
  reg [31:0] _T_422_im; // @[Reg.scala 15:16]
  reg [31:0] _T_423_re; // @[Reg.scala 15:16]
  reg [31:0] _T_423_im; // @[Reg.scala 15:16]
  reg [31:0] _T_424_re; // @[Reg.scala 15:16]
  reg [31:0] _T_424_im; // @[Reg.scala 15:16]
  reg [31:0] _T_425_re; // @[Reg.scala 15:16]
  reg [31:0] _T_425_im; // @[Reg.scala 15:16]
  reg [31:0] _T_426_re; // @[Reg.scala 15:16]
  reg [31:0] _T_426_im; // @[Reg.scala 15:16]
  reg [31:0] _T_427_re; // @[Reg.scala 15:16]
  reg [31:0] _T_427_im; // @[Reg.scala 15:16]
  reg [31:0] _T_428_re; // @[Reg.scala 15:16]
  reg [31:0] _T_428_im; // @[Reg.scala 15:16]
  reg [31:0] _T_429_re; // @[Reg.scala 15:16]
  reg [31:0] _T_429_im; // @[Reg.scala 15:16]
  reg [31:0] _T_430_re; // @[Reg.scala 15:16]
  reg [31:0] _T_430_im; // @[Reg.scala 15:16]
  reg [31:0] _T_431_re; // @[Reg.scala 15:16]
  reg [31:0] _T_431_im; // @[Reg.scala 15:16]
  reg [31:0] _T_432_re; // @[Reg.scala 15:16]
  reg [31:0] _T_432_im; // @[Reg.scala 15:16]
  reg [31:0] _T_433_re; // @[Reg.scala 15:16]
  reg [31:0] _T_433_im; // @[Reg.scala 15:16]
  reg [31:0] _T_434_re; // @[Reg.scala 15:16]
  reg [31:0] _T_434_im; // @[Reg.scala 15:16]
  reg [31:0] _T_435_re; // @[Reg.scala 15:16]
  reg [31:0] _T_435_im; // @[Reg.scala 15:16]
  reg [31:0] _T_436_re; // @[Reg.scala 15:16]
  reg [31:0] _T_436_im; // @[Reg.scala 15:16]
  reg [31:0] _T_437_re; // @[Reg.scala 15:16]
  reg [31:0] _T_437_im; // @[Reg.scala 15:16]
  reg [31:0] _T_438_re; // @[Reg.scala 15:16]
  reg [31:0] _T_438_im; // @[Reg.scala 15:16]
  reg [31:0] _T_439_re; // @[Reg.scala 15:16]
  reg [31:0] _T_439_im; // @[Reg.scala 15:16]
  reg [31:0] _T_440_re; // @[Reg.scala 15:16]
  reg [31:0] _T_440_im; // @[Reg.scala 15:16]
  reg [31:0] _T_441_re; // @[Reg.scala 15:16]
  reg [31:0] _T_441_im; // @[Reg.scala 15:16]
  reg [31:0] _T_442_re; // @[Reg.scala 15:16]
  reg [31:0] _T_442_im; // @[Reg.scala 15:16]
  reg [31:0] _T_443_re; // @[Reg.scala 15:16]
  reg [31:0] _T_443_im; // @[Reg.scala 15:16]
  reg [31:0] _T_444_re; // @[Reg.scala 15:16]
  reg [31:0] _T_444_im; // @[Reg.scala 15:16]
  reg [31:0] _T_445_re; // @[Reg.scala 15:16]
  reg [31:0] _T_445_im; // @[Reg.scala 15:16]
  reg [31:0] _T_446_re; // @[Reg.scala 15:16]
  reg [31:0] _T_446_im; // @[Reg.scala 15:16]
  reg [31:0] _T_447_re; // @[Reg.scala 15:16]
  reg [31:0] _T_447_im; // @[Reg.scala 15:16]
  reg [31:0] _T_448_re; // @[Reg.scala 15:16]
  reg [31:0] _T_448_im; // @[Reg.scala 15:16]
  reg [31:0] _T_449_re; // @[Reg.scala 15:16]
  reg [31:0] _T_449_im; // @[Reg.scala 15:16]
  reg [31:0] _T_450_re; // @[Reg.scala 15:16]
  reg [31:0] _T_450_im; // @[Reg.scala 15:16]
  reg [31:0] _T_451_re; // @[Reg.scala 15:16]
  reg [31:0] _T_451_im; // @[Reg.scala 15:16]
  reg [31:0] _T_452_re; // @[Reg.scala 15:16]
  reg [31:0] _T_452_im; // @[Reg.scala 15:16]
  reg [31:0] _T_453_re; // @[Reg.scala 15:16]
  reg [31:0] _T_453_im; // @[Reg.scala 15:16]
  reg [31:0] _T_454_re; // @[Reg.scala 15:16]
  reg [31:0] _T_454_im; // @[Reg.scala 15:16]
  reg [31:0] _T_455_re; // @[Reg.scala 15:16]
  reg [31:0] _T_455_im; // @[Reg.scala 15:16]
  reg [31:0] _T_456_re; // @[Reg.scala 15:16]
  reg [31:0] _T_456_im; // @[Reg.scala 15:16]
  reg [31:0] _T_457_re; // @[Reg.scala 15:16]
  reg [31:0] _T_457_im; // @[Reg.scala 15:16]
  reg [31:0] _T_458_re; // @[Reg.scala 15:16]
  reg [31:0] _T_458_im; // @[Reg.scala 15:16]
  reg [31:0] _T_459_re; // @[Reg.scala 15:16]
  reg [31:0] _T_459_im; // @[Reg.scala 15:16]
  reg [31:0] _T_460_re; // @[Reg.scala 15:16]
  reg [31:0] _T_460_im; // @[Reg.scala 15:16]
  reg [31:0] _T_461_re; // @[Reg.scala 15:16]
  reg [31:0] _T_461_im; // @[Reg.scala 15:16]
  reg [31:0] _T_462_re; // @[Reg.scala 15:16]
  reg [31:0] _T_462_im; // @[Reg.scala 15:16]
  reg [31:0] _T_463_re; // @[Reg.scala 15:16]
  reg [31:0] _T_463_im; // @[Reg.scala 15:16]
  reg [31:0] _T_464_re; // @[Reg.scala 15:16]
  reg [31:0] _T_464_im; // @[Reg.scala 15:16]
  reg [31:0] _T_465_re; // @[Reg.scala 15:16]
  reg [31:0] _T_465_im; // @[Reg.scala 15:16]
  reg [31:0] _T_466_re; // @[Reg.scala 15:16]
  reg [31:0] _T_466_im; // @[Reg.scala 15:16]
  reg [31:0] _T_467_re; // @[Reg.scala 15:16]
  reg [31:0] _T_467_im; // @[Reg.scala 15:16]
  reg [31:0] _T_468_re; // @[Reg.scala 15:16]
  reg [31:0] _T_468_im; // @[Reg.scala 15:16]
  reg [31:0] _T_469_re; // @[Reg.scala 15:16]
  reg [31:0] _T_469_im; // @[Reg.scala 15:16]
  reg [31:0] _T_470_re; // @[Reg.scala 15:16]
  reg [31:0] _T_470_im; // @[Reg.scala 15:16]
  reg [31:0] _T_471_re; // @[Reg.scala 15:16]
  reg [31:0] _T_471_im; // @[Reg.scala 15:16]
  reg [31:0] _T_472_re; // @[Reg.scala 15:16]
  reg [31:0] _T_472_im; // @[Reg.scala 15:16]
  reg [31:0] _T_473_re; // @[Reg.scala 15:16]
  reg [31:0] _T_473_im; // @[Reg.scala 15:16]
  reg [31:0] _T_474_re; // @[Reg.scala 15:16]
  reg [31:0] _T_474_im; // @[Reg.scala 15:16]
  reg [31:0] _T_475_re; // @[Reg.scala 15:16]
  reg [31:0] _T_475_im; // @[Reg.scala 15:16]
  reg [31:0] _T_476_re; // @[Reg.scala 15:16]
  reg [31:0] _T_476_im; // @[Reg.scala 15:16]
  reg [31:0] _T_477_re; // @[Reg.scala 15:16]
  reg [31:0] _T_477_im; // @[Reg.scala 15:16]
  reg [31:0] _T_478_re; // @[Reg.scala 15:16]
  reg [31:0] _T_478_im; // @[Reg.scala 15:16]
  reg [31:0] _T_479_re; // @[Reg.scala 15:16]
  reg [31:0] _T_479_im; // @[Reg.scala 15:16]
  reg [31:0] _T_480_re; // @[Reg.scala 15:16]
  reg [31:0] _T_480_im; // @[Reg.scala 15:16]
  reg [31:0] _T_481_re; // @[Reg.scala 15:16]
  reg [31:0] _T_481_im; // @[Reg.scala 15:16]
  reg [31:0] _T_482_re; // @[Reg.scala 15:16]
  reg [31:0] _T_482_im; // @[Reg.scala 15:16]
  reg [31:0] _T_483_re; // @[Reg.scala 15:16]
  reg [31:0] _T_483_im; // @[Reg.scala 15:16]
  reg [31:0] _T_484_re; // @[Reg.scala 15:16]
  reg [31:0] _T_484_im; // @[Reg.scala 15:16]
  reg [31:0] _T_485_re; // @[Reg.scala 15:16]
  reg [31:0] _T_485_im; // @[Reg.scala 15:16]
  reg [31:0] _T_486_re; // @[Reg.scala 15:16]
  reg [31:0] _T_486_im; // @[Reg.scala 15:16]
  reg [31:0] _T_487_re; // @[Reg.scala 15:16]
  reg [31:0] _T_487_im; // @[Reg.scala 15:16]
  reg [31:0] _T_488_re; // @[Reg.scala 15:16]
  reg [31:0] _T_488_im; // @[Reg.scala 15:16]
  reg [31:0] _T_489_re; // @[Reg.scala 15:16]
  reg [31:0] _T_489_im; // @[Reg.scala 15:16]
  reg [31:0] _T_490_re; // @[Reg.scala 15:16]
  reg [31:0] _T_490_im; // @[Reg.scala 15:16]
  reg [31:0] _T_491_re; // @[Reg.scala 15:16]
  reg [31:0] _T_491_im; // @[Reg.scala 15:16]
  reg [31:0] _T_492_re; // @[Reg.scala 15:16]
  reg [31:0] _T_492_im; // @[Reg.scala 15:16]
  reg [31:0] _T_493_re; // @[Reg.scala 15:16]
  reg [31:0] _T_493_im; // @[Reg.scala 15:16]
  reg [31:0] _T_494_re; // @[Reg.scala 15:16]
  reg [31:0] _T_494_im; // @[Reg.scala 15:16]
  reg [31:0] _T_495_re; // @[Reg.scala 15:16]
  reg [31:0] _T_495_im; // @[Reg.scala 15:16]
  reg [31:0] _T_496_re; // @[Reg.scala 15:16]
  reg [31:0] _T_496_im; // @[Reg.scala 15:16]
  reg [31:0] _T_497_re; // @[Reg.scala 15:16]
  reg [31:0] _T_497_im; // @[Reg.scala 15:16]
  reg [31:0] _T_498_re; // @[Reg.scala 15:16]
  reg [31:0] _T_498_im; // @[Reg.scala 15:16]
  reg [31:0] _T_499_re; // @[Reg.scala 15:16]
  reg [31:0] _T_499_im; // @[Reg.scala 15:16]
  reg [31:0] _T_500_re; // @[Reg.scala 15:16]
  reg [31:0] _T_500_im; // @[Reg.scala 15:16]
  reg [31:0] _T_501_re; // @[Reg.scala 15:16]
  reg [31:0] _T_501_im; // @[Reg.scala 15:16]
  reg [31:0] _T_502_re; // @[Reg.scala 15:16]
  reg [31:0] _T_502_im; // @[Reg.scala 15:16]
  reg [31:0] _T_503_re; // @[Reg.scala 15:16]
  reg [31:0] _T_503_im; // @[Reg.scala 15:16]
  reg [31:0] _T_504_re; // @[Reg.scala 15:16]
  reg [31:0] _T_504_im; // @[Reg.scala 15:16]
  reg [31:0] _T_505_re; // @[Reg.scala 15:16]
  reg [31:0] _T_505_im; // @[Reg.scala 15:16]
  reg [31:0] _T_506_re; // @[Reg.scala 15:16]
  reg [31:0] _T_506_im; // @[Reg.scala 15:16]
  reg [31:0] _T_507_re; // @[Reg.scala 15:16]
  reg [31:0] _T_507_im; // @[Reg.scala 15:16]
  reg [31:0] _T_508_re; // @[Reg.scala 15:16]
  reg [31:0] _T_508_im; // @[Reg.scala 15:16]
  reg [31:0] _T_509_re; // @[Reg.scala 15:16]
  reg [31:0] _T_509_im; // @[Reg.scala 15:16]
  reg [31:0] _T_510_re; // @[Reg.scala 15:16]
  reg [31:0] _T_510_im; // @[Reg.scala 15:16]
  reg [31:0] _T_511_re; // @[Reg.scala 15:16]
  reg [31:0] _T_511_im; // @[Reg.scala 15:16]
  reg [31:0] _T_512_re; // @[Reg.scala 15:16]
  reg [31:0] _T_512_im; // @[Reg.scala 15:16]
  reg [31:0] _T_513_re; // @[Reg.scala 15:16]
  reg [31:0] _T_513_im; // @[Reg.scala 15:16]
  reg [31:0] _T_514_re; // @[Reg.scala 15:16]
  reg [31:0] _T_514_im; // @[Reg.scala 15:16]
  reg [31:0] _T_515_re; // @[Reg.scala 15:16]
  reg [31:0] _T_515_im; // @[Reg.scala 15:16]
  reg [31:0] _T_516_re; // @[Reg.scala 15:16]
  reg [31:0] _T_516_im; // @[Reg.scala 15:16]
  reg [31:0] _T_517_re; // @[Reg.scala 15:16]
  reg [31:0] _T_517_im; // @[Reg.scala 15:16]
  reg [31:0] _T_518_re; // @[Reg.scala 15:16]
  reg [31:0] _T_518_im; // @[Reg.scala 15:16]
  reg [31:0] _T_519_re; // @[Reg.scala 15:16]
  reg [31:0] _T_519_im; // @[Reg.scala 15:16]
  reg [31:0] _T_520_re; // @[Reg.scala 15:16]
  reg [31:0] _T_520_im; // @[Reg.scala 15:16]
  reg [31:0] _T_521_re; // @[Reg.scala 15:16]
  reg [31:0] _T_521_im; // @[Reg.scala 15:16]
  reg [31:0] _T_522_re; // @[Reg.scala 15:16]
  reg [31:0] _T_522_im; // @[Reg.scala 15:16]
  reg [31:0] _T_523_re; // @[Reg.scala 15:16]
  reg [31:0] _T_523_im; // @[Reg.scala 15:16]
  reg [31:0] _T_524_re; // @[Reg.scala 15:16]
  reg [31:0] _T_524_im; // @[Reg.scala 15:16]
  reg [31:0] _T_525_re; // @[Reg.scala 15:16]
  reg [31:0] _T_525_im; // @[Reg.scala 15:16]
  reg [31:0] _T_526_re; // @[Reg.scala 15:16]
  reg [31:0] _T_526_im; // @[Reg.scala 15:16]
  reg [31:0] _T_527_re; // @[Reg.scala 15:16]
  reg [31:0] _T_527_im; // @[Reg.scala 15:16]
  reg [31:0] _T_528_re; // @[Reg.scala 15:16]
  reg [31:0] _T_528_im; // @[Reg.scala 15:16]
  reg [31:0] _T_529_re; // @[Reg.scala 15:16]
  reg [31:0] _T_529_im; // @[Reg.scala 15:16]
  reg [31:0] _T_530_re; // @[Reg.scala 15:16]
  reg [31:0] _T_530_im; // @[Reg.scala 15:16]
  reg [31:0] _T_531_re; // @[Reg.scala 15:16]
  reg [31:0] _T_531_im; // @[Reg.scala 15:16]
  reg [31:0] _T_532_re; // @[Reg.scala 15:16]
  reg [31:0] _T_532_im; // @[Reg.scala 15:16]
  reg [31:0] _T_533_re; // @[Reg.scala 15:16]
  reg [31:0] _T_533_im; // @[Reg.scala 15:16]
  reg [31:0] _T_534_re; // @[Reg.scala 15:16]
  reg [31:0] _T_534_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_1794 = 7'h1 == cnt[6:0] ? $signed(32'shffec) : $signed(32'sh10000); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1795 = 7'h2 == cnt[6:0] ? $signed(32'shffb1) : $signed(_GEN_1794); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1796 = 7'h3 == cnt[6:0] ? $signed(32'shff4e) : $signed(_GEN_1795); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1797 = 7'h4 == cnt[6:0] ? $signed(32'shfec4) : $signed(_GEN_1796); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1798 = 7'h5 == cnt[6:0] ? $signed(32'shfe13) : $signed(_GEN_1797); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1799 = 7'h6 == cnt[6:0] ? $signed(32'shfd3b) : $signed(_GEN_1798); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1800 = 7'h7 == cnt[6:0] ? $signed(32'shfc3b) : $signed(_GEN_1799); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1801 = 7'h8 == cnt[6:0] ? $signed(32'shfb15) : $signed(_GEN_1800); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1802 = 7'h9 == cnt[6:0] ? $signed(32'shf9c8) : $signed(_GEN_1801); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1803 = 7'ha == cnt[6:0] ? $signed(32'shf854) : $signed(_GEN_1802); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1804 = 7'hb == cnt[6:0] ? $signed(32'shf6ba) : $signed(_GEN_1803); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1805 = 7'hc == cnt[6:0] ? $signed(32'shf4fa) : $signed(_GEN_1804); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1806 = 7'hd == cnt[6:0] ? $signed(32'shf314) : $signed(_GEN_1805); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1807 = 7'he == cnt[6:0] ? $signed(32'shf109) : $signed(_GEN_1806); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1808 = 7'hf == cnt[6:0] ? $signed(32'sheed9) : $signed(_GEN_1807); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1809 = 7'h10 == cnt[6:0] ? $signed(32'shec83) : $signed(_GEN_1808); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1810 = 7'h11 == cnt[6:0] ? $signed(32'shea0a) : $signed(_GEN_1809); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1811 = 7'h12 == cnt[6:0] ? $signed(32'she76c) : $signed(_GEN_1810); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1812 = 7'h13 == cnt[6:0] ? $signed(32'she4aa) : $signed(_GEN_1811); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1813 = 7'h14 == cnt[6:0] ? $signed(32'she1c6) : $signed(_GEN_1812); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1814 = 7'h15 == cnt[6:0] ? $signed(32'shdebe) : $signed(_GEN_1813); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1815 = 7'h16 == cnt[6:0] ? $signed(32'shdb94) : $signed(_GEN_1814); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1816 = 7'h17 == cnt[6:0] ? $signed(32'shd848) : $signed(_GEN_1815); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1817 = 7'h18 == cnt[6:0] ? $signed(32'shd4db) : $signed(_GEN_1816); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1818 = 7'h19 == cnt[6:0] ? $signed(32'shd14d) : $signed(_GEN_1817); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1819 = 7'h1a == cnt[6:0] ? $signed(32'shcd9f) : $signed(_GEN_1818); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1820 = 7'h1b == cnt[6:0] ? $signed(32'shc9d1) : $signed(_GEN_1819); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1821 = 7'h1c == cnt[6:0] ? $signed(32'shc5e4) : $signed(_GEN_1820); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1822 = 7'h1d == cnt[6:0] ? $signed(32'shc1d8) : $signed(_GEN_1821); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1823 = 7'h1e == cnt[6:0] ? $signed(32'shbdaf) : $signed(_GEN_1822); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1824 = 7'h1f == cnt[6:0] ? $signed(32'shb968) : $signed(_GEN_1823); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1825 = 7'h20 == cnt[6:0] ? $signed(32'shb505) : $signed(_GEN_1824); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1826 = 7'h21 == cnt[6:0] ? $signed(32'shb086) : $signed(_GEN_1825); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1827 = 7'h22 == cnt[6:0] ? $signed(32'shabeb) : $signed(_GEN_1826); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1828 = 7'h23 == cnt[6:0] ? $signed(32'sha736) : $signed(_GEN_1827); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1829 = 7'h24 == cnt[6:0] ? $signed(32'sha268) : $signed(_GEN_1828); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1830 = 7'h25 == cnt[6:0] ? $signed(32'sh9d80) : $signed(_GEN_1829); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1831 = 7'h26 == cnt[6:0] ? $signed(32'sh9880) : $signed(_GEN_1830); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1832 = 7'h27 == cnt[6:0] ? $signed(32'sh9368) : $signed(_GEN_1831); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1833 = 7'h28 == cnt[6:0] ? $signed(32'sh8e3a) : $signed(_GEN_1832); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1834 = 7'h29 == cnt[6:0] ? $signed(32'sh88f6) : $signed(_GEN_1833); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1835 = 7'h2a == cnt[6:0] ? $signed(32'sh839c) : $signed(_GEN_1834); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1836 = 7'h2b == cnt[6:0] ? $signed(32'sh7e2f) : $signed(_GEN_1835); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1837 = 7'h2c == cnt[6:0] ? $signed(32'sh78ad) : $signed(_GEN_1836); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1838 = 7'h2d == cnt[6:0] ? $signed(32'sh731a) : $signed(_GEN_1837); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1839 = 7'h2e == cnt[6:0] ? $signed(32'sh6d74) : $signed(_GEN_1838); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1840 = 7'h2f == cnt[6:0] ? $signed(32'sh67be) : $signed(_GEN_1839); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1841 = 7'h30 == cnt[6:0] ? $signed(32'sh61f8) : $signed(_GEN_1840); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1842 = 7'h31 == cnt[6:0] ? $signed(32'sh5c22) : $signed(_GEN_1841); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1843 = 7'h32 == cnt[6:0] ? $signed(32'sh563e) : $signed(_GEN_1842); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1844 = 7'h33 == cnt[6:0] ? $signed(32'sh504d) : $signed(_GEN_1843); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1845 = 7'h34 == cnt[6:0] ? $signed(32'sh4a50) : $signed(_GEN_1844); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1846 = 7'h35 == cnt[6:0] ? $signed(32'sh4447) : $signed(_GEN_1845); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1847 = 7'h36 == cnt[6:0] ? $signed(32'sh3e34) : $signed(_GEN_1846); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1848 = 7'h37 == cnt[6:0] ? $signed(32'sh3817) : $signed(_GEN_1847); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1849 = 7'h38 == cnt[6:0] ? $signed(32'sh31f1) : $signed(_GEN_1848); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1850 = 7'h39 == cnt[6:0] ? $signed(32'sh2bc4) : $signed(_GEN_1849); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1851 = 7'h3a == cnt[6:0] ? $signed(32'sh2590) : $signed(_GEN_1850); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1852 = 7'h3b == cnt[6:0] ? $signed(32'sh1f56) : $signed(_GEN_1851); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1853 = 7'h3c == cnt[6:0] ? $signed(32'sh1918) : $signed(_GEN_1852); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1854 = 7'h3d == cnt[6:0] ? $signed(32'sh12d5) : $signed(_GEN_1853); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1855 = 7'h3e == cnt[6:0] ? $signed(32'shc90) : $signed(_GEN_1854); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1856 = 7'h3f == cnt[6:0] ? $signed(32'sh648) : $signed(_GEN_1855); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1857 = 7'h40 == cnt[6:0] ? $signed(32'sh0) : $signed(_GEN_1856); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1858 = 7'h41 == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_1857); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1859 = 7'h42 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_1858); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1860 = 7'h43 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_1859); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1861 = 7'h44 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_1860); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1862 = 7'h45 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_1861); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1863 = 7'h46 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_1862); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1864 = 7'h47 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_1863); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1865 = 7'h48 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_1864); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1866 = 7'h49 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_1865); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1867 = 7'h4a == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_1866); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1868 = 7'h4b == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_1867); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1869 = 7'h4c == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_1868); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1870 = 7'h4d == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_1869); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1871 = 7'h4e == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_1870); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1872 = 7'h4f == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_1871); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1873 = 7'h50 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_1872); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1874 = 7'h51 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_1873); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1875 = 7'h52 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_1874); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1876 = 7'h53 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_1875); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1877 = 7'h54 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_1876); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1878 = 7'h55 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_1877); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1879 = 7'h56 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_1878); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1880 = 7'h57 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_1879); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1881 = 7'h58 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_1880); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1882 = 7'h59 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_1881); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1883 = 7'h5a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_1882); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1884 = 7'h5b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_1883); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1885 = 7'h5c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_1884); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1886 = 7'h5d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_1885); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1887 = 7'h5e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_1886); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1888 = 7'h5f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_1887); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1889 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_1888); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1890 = 7'h61 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_1889); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1891 = 7'h62 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_1890); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1892 = 7'h63 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_1891); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1893 = 7'h64 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_1892); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1894 = 7'h65 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_1893); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1895 = 7'h66 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_1894); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1896 = 7'h67 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_1895); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1897 = 7'h68 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_1896); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1898 = 7'h69 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_1897); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1899 = 7'h6a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_1898); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1900 = 7'h6b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_1899); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1901 = 7'h6c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_1900); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1902 = 7'h6d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_1901); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1903 = 7'h6e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_1902); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1904 = 7'h6f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_1903); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1905 = 7'h70 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_1904); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1906 = 7'h71 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_1905); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1907 = 7'h72 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_1906); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1908 = 7'h73 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_1907); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1909 = 7'h74 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_1908); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1910 = 7'h75 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_1909); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1911 = 7'h76 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_1910); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1912 = 7'h77 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_1911); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1913 = 7'h78 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_1912); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1914 = 7'h79 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_1913); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1915 = 7'h7a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_1914); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1916 = 7'h7b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_1915); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1917 = 7'h7c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_1916); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1918 = 7'h7d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_1917); // @[FFT.scala 51:18]
  wire [31:0] _GEN_1919 = 7'h7e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_1918); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2178 = 7'h1 == cnt[6:0] ? $signed(-32'sh648) : $signed(32'sh0); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2179 = 7'h2 == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_2178); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2180 = 7'h3 == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_2179); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2181 = 7'h4 == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_2180); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2182 = 7'h5 == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_2181); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2183 = 7'h6 == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_2182); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2184 = 7'h7 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_2183); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2185 = 7'h8 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_2184); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2186 = 7'h9 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_2185); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2187 = 7'ha == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_2186); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2188 = 7'hb == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_2187); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2189 = 7'hc == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_2188); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2190 = 7'hd == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_2189); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2191 = 7'he == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_2190); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2192 = 7'hf == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_2191); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2193 = 7'h10 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_2192); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2194 = 7'h11 == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_2193); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2195 = 7'h12 == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_2194); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2196 = 7'h13 == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_2195); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2197 = 7'h14 == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_2196); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2198 = 7'h15 == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_2197); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2199 = 7'h16 == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_2198); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2200 = 7'h17 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_2199); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2201 = 7'h18 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2200); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2202 = 7'h19 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_2201); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2203 = 7'h1a == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_2202); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2204 = 7'h1b == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_2203); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2205 = 7'h1c == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_2204); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2206 = 7'h1d == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_2205); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2207 = 7'h1e == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_2206); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2208 = 7'h1f == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_2207); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2209 = 7'h20 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_2208); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2210 = 7'h21 == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_2209); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2211 = 7'h22 == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_2210); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2212 = 7'h23 == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_2211); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2213 = 7'h24 == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_2212); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2214 = 7'h25 == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_2213); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2215 = 7'h26 == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_2214); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2216 = 7'h27 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_2215); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2217 = 7'h28 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_2216); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2218 = 7'h29 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_2217); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2219 = 7'h2a == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_2218); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2220 = 7'h2b == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_2219); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2221 = 7'h2c == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_2220); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2222 = 7'h2d == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_2221); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2223 = 7'h2e == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_2222); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2224 = 7'h2f == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_2223); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2225 = 7'h30 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_2224); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2226 = 7'h31 == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_2225); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2227 = 7'h32 == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_2226); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2228 = 7'h33 == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_2227); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2229 = 7'h34 == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_2228); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2230 = 7'h35 == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_2229); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2231 = 7'h36 == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_2230); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2232 = 7'h37 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_2231); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2233 = 7'h38 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_2232); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2234 = 7'h39 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_2233); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2235 = 7'h3a == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_2234); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2236 = 7'h3b == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_2235); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2237 = 7'h3c == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_2236); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2238 = 7'h3d == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_2237); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2239 = 7'h3e == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_2238); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2240 = 7'h3f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_2239); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2241 = 7'h40 == cnt[6:0] ? $signed(-32'sh10000) : $signed(_GEN_2240); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2242 = 7'h41 == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_2241); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2243 = 7'h42 == cnt[6:0] ? $signed(-32'shffb1) : $signed(_GEN_2242); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2244 = 7'h43 == cnt[6:0] ? $signed(-32'shff4e) : $signed(_GEN_2243); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2245 = 7'h44 == cnt[6:0] ? $signed(-32'shfec4) : $signed(_GEN_2244); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2246 = 7'h45 == cnt[6:0] ? $signed(-32'shfe13) : $signed(_GEN_2245); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2247 = 7'h46 == cnt[6:0] ? $signed(-32'shfd3b) : $signed(_GEN_2246); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2248 = 7'h47 == cnt[6:0] ? $signed(-32'shfc3b) : $signed(_GEN_2247); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2249 = 7'h48 == cnt[6:0] ? $signed(-32'shfb15) : $signed(_GEN_2248); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2250 = 7'h49 == cnt[6:0] ? $signed(-32'shf9c8) : $signed(_GEN_2249); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2251 = 7'h4a == cnt[6:0] ? $signed(-32'shf854) : $signed(_GEN_2250); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2252 = 7'h4b == cnt[6:0] ? $signed(-32'shf6ba) : $signed(_GEN_2251); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2253 = 7'h4c == cnt[6:0] ? $signed(-32'shf4fa) : $signed(_GEN_2252); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2254 = 7'h4d == cnt[6:0] ? $signed(-32'shf314) : $signed(_GEN_2253); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2255 = 7'h4e == cnt[6:0] ? $signed(-32'shf109) : $signed(_GEN_2254); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2256 = 7'h4f == cnt[6:0] ? $signed(-32'sheed9) : $signed(_GEN_2255); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2257 = 7'h50 == cnt[6:0] ? $signed(-32'shec83) : $signed(_GEN_2256); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2258 = 7'h51 == cnt[6:0] ? $signed(-32'shea0a) : $signed(_GEN_2257); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2259 = 7'h52 == cnt[6:0] ? $signed(-32'she76c) : $signed(_GEN_2258); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2260 = 7'h53 == cnt[6:0] ? $signed(-32'she4aa) : $signed(_GEN_2259); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2261 = 7'h54 == cnt[6:0] ? $signed(-32'she1c6) : $signed(_GEN_2260); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2262 = 7'h55 == cnt[6:0] ? $signed(-32'shdebe) : $signed(_GEN_2261); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2263 = 7'h56 == cnt[6:0] ? $signed(-32'shdb94) : $signed(_GEN_2262); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2264 = 7'h57 == cnt[6:0] ? $signed(-32'shd848) : $signed(_GEN_2263); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2265 = 7'h58 == cnt[6:0] ? $signed(-32'shd4db) : $signed(_GEN_2264); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2266 = 7'h59 == cnt[6:0] ? $signed(-32'shd14d) : $signed(_GEN_2265); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2267 = 7'h5a == cnt[6:0] ? $signed(-32'shcd9f) : $signed(_GEN_2266); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2268 = 7'h5b == cnt[6:0] ? $signed(-32'shc9d1) : $signed(_GEN_2267); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2269 = 7'h5c == cnt[6:0] ? $signed(-32'shc5e4) : $signed(_GEN_2268); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2270 = 7'h5d == cnt[6:0] ? $signed(-32'shc1d8) : $signed(_GEN_2269); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2271 = 7'h5e == cnt[6:0] ? $signed(-32'shbdaf) : $signed(_GEN_2270); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2272 = 7'h5f == cnt[6:0] ? $signed(-32'shb968) : $signed(_GEN_2271); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2273 = 7'h60 == cnt[6:0] ? $signed(-32'shb505) : $signed(_GEN_2272); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2274 = 7'h61 == cnt[6:0] ? $signed(-32'shb086) : $signed(_GEN_2273); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2275 = 7'h62 == cnt[6:0] ? $signed(-32'shabeb) : $signed(_GEN_2274); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2276 = 7'h63 == cnt[6:0] ? $signed(-32'sha736) : $signed(_GEN_2275); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2277 = 7'h64 == cnt[6:0] ? $signed(-32'sha268) : $signed(_GEN_2276); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2278 = 7'h65 == cnt[6:0] ? $signed(-32'sh9d80) : $signed(_GEN_2277); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2279 = 7'h66 == cnt[6:0] ? $signed(-32'sh9880) : $signed(_GEN_2278); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2280 = 7'h67 == cnt[6:0] ? $signed(-32'sh9368) : $signed(_GEN_2279); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2281 = 7'h68 == cnt[6:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2280); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2282 = 7'h69 == cnt[6:0] ? $signed(-32'sh88f6) : $signed(_GEN_2281); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2283 = 7'h6a == cnt[6:0] ? $signed(-32'sh839c) : $signed(_GEN_2282); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2284 = 7'h6b == cnt[6:0] ? $signed(-32'sh7e2f) : $signed(_GEN_2283); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2285 = 7'h6c == cnt[6:0] ? $signed(-32'sh78ad) : $signed(_GEN_2284); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2286 = 7'h6d == cnt[6:0] ? $signed(-32'sh731a) : $signed(_GEN_2285); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2287 = 7'h6e == cnt[6:0] ? $signed(-32'sh6d74) : $signed(_GEN_2286); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2288 = 7'h6f == cnt[6:0] ? $signed(-32'sh67be) : $signed(_GEN_2287); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2289 = 7'h70 == cnt[6:0] ? $signed(-32'sh61f8) : $signed(_GEN_2288); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2290 = 7'h71 == cnt[6:0] ? $signed(-32'sh5c22) : $signed(_GEN_2289); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2291 = 7'h72 == cnt[6:0] ? $signed(-32'sh563e) : $signed(_GEN_2290); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2292 = 7'h73 == cnt[6:0] ? $signed(-32'sh504d) : $signed(_GEN_2291); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2293 = 7'h74 == cnt[6:0] ? $signed(-32'sh4a50) : $signed(_GEN_2292); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2294 = 7'h75 == cnt[6:0] ? $signed(-32'sh4447) : $signed(_GEN_2293); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2295 = 7'h76 == cnt[6:0] ? $signed(-32'sh3e34) : $signed(_GEN_2294); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2296 = 7'h77 == cnt[6:0] ? $signed(-32'sh3817) : $signed(_GEN_2295); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2297 = 7'h78 == cnt[6:0] ? $signed(-32'sh31f1) : $signed(_GEN_2296); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2298 = 7'h79 == cnt[6:0] ? $signed(-32'sh2bc4) : $signed(_GEN_2297); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2299 = 7'h7a == cnt[6:0] ? $signed(-32'sh2590) : $signed(_GEN_2298); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2300 = 7'h7b == cnt[6:0] ? $signed(-32'sh1f56) : $signed(_GEN_2299); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2301 = 7'h7c == cnt[6:0] ? $signed(-32'sh1918) : $signed(_GEN_2300); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2302 = 7'h7d == cnt[6:0] ? $signed(-32'sh12d5) : $signed(_GEN_2301); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2303 = 7'h7e == cnt[6:0] ? $signed(-32'shc90) : $signed(_GEN_2302); // @[FFT.scala 52:18]
  reg [31:0] _T_543_re; // @[Reg.scala 15:16]
  reg [31:0] _T_543_im; // @[Reg.scala 15:16]
  reg [31:0] _T_544_re; // @[Reg.scala 15:16]
  reg [31:0] _T_544_im; // @[Reg.scala 15:16]
  reg [31:0] _T_545_re; // @[Reg.scala 15:16]
  reg [31:0] _T_545_im; // @[Reg.scala 15:16]
  reg [31:0] _T_546_re; // @[Reg.scala 15:16]
  reg [31:0] _T_546_im; // @[Reg.scala 15:16]
  reg [31:0] _T_547_re; // @[Reg.scala 15:16]
  reg [31:0] _T_547_im; // @[Reg.scala 15:16]
  reg [31:0] _T_548_re; // @[Reg.scala 15:16]
  reg [31:0] _T_548_im; // @[Reg.scala 15:16]
  reg [31:0] _T_549_re; // @[Reg.scala 15:16]
  reg [31:0] _T_549_im; // @[Reg.scala 15:16]
  reg [31:0] _T_550_re; // @[Reg.scala 15:16]
  reg [31:0] _T_550_im; // @[Reg.scala 15:16]
  reg [31:0] _T_551_re; // @[Reg.scala 15:16]
  reg [31:0] _T_551_im; // @[Reg.scala 15:16]
  reg [31:0] _T_552_re; // @[Reg.scala 15:16]
  reg [31:0] _T_552_im; // @[Reg.scala 15:16]
  reg [31:0] _T_553_re; // @[Reg.scala 15:16]
  reg [31:0] _T_553_im; // @[Reg.scala 15:16]
  reg [31:0] _T_554_re; // @[Reg.scala 15:16]
  reg [31:0] _T_554_im; // @[Reg.scala 15:16]
  reg [31:0] _T_555_re; // @[Reg.scala 15:16]
  reg [31:0] _T_555_im; // @[Reg.scala 15:16]
  reg [31:0] _T_556_re; // @[Reg.scala 15:16]
  reg [31:0] _T_556_im; // @[Reg.scala 15:16]
  reg [31:0] _T_557_re; // @[Reg.scala 15:16]
  reg [31:0] _T_557_im; // @[Reg.scala 15:16]
  reg [31:0] _T_558_re; // @[Reg.scala 15:16]
  reg [31:0] _T_558_im; // @[Reg.scala 15:16]
  reg [31:0] _T_559_re; // @[Reg.scala 15:16]
  reg [31:0] _T_559_im; // @[Reg.scala 15:16]
  reg [31:0] _T_560_re; // @[Reg.scala 15:16]
  reg [31:0] _T_560_im; // @[Reg.scala 15:16]
  reg [31:0] _T_561_re; // @[Reg.scala 15:16]
  reg [31:0] _T_561_im; // @[Reg.scala 15:16]
  reg [31:0] _T_562_re; // @[Reg.scala 15:16]
  reg [31:0] _T_562_im; // @[Reg.scala 15:16]
  reg [31:0] _T_563_re; // @[Reg.scala 15:16]
  reg [31:0] _T_563_im; // @[Reg.scala 15:16]
  reg [31:0] _T_564_re; // @[Reg.scala 15:16]
  reg [31:0] _T_564_im; // @[Reg.scala 15:16]
  reg [31:0] _T_565_re; // @[Reg.scala 15:16]
  reg [31:0] _T_565_im; // @[Reg.scala 15:16]
  reg [31:0] _T_566_re; // @[Reg.scala 15:16]
  reg [31:0] _T_566_im; // @[Reg.scala 15:16]
  reg [31:0] _T_567_re; // @[Reg.scala 15:16]
  reg [31:0] _T_567_im; // @[Reg.scala 15:16]
  reg [31:0] _T_568_re; // @[Reg.scala 15:16]
  reg [31:0] _T_568_im; // @[Reg.scala 15:16]
  reg [31:0] _T_569_re; // @[Reg.scala 15:16]
  reg [31:0] _T_569_im; // @[Reg.scala 15:16]
  reg [31:0] _T_570_re; // @[Reg.scala 15:16]
  reg [31:0] _T_570_im; // @[Reg.scala 15:16]
  reg [31:0] _T_571_re; // @[Reg.scala 15:16]
  reg [31:0] _T_571_im; // @[Reg.scala 15:16]
  reg [31:0] _T_572_re; // @[Reg.scala 15:16]
  reg [31:0] _T_572_im; // @[Reg.scala 15:16]
  reg [31:0] _T_573_re; // @[Reg.scala 15:16]
  reg [31:0] _T_573_im; // @[Reg.scala 15:16]
  reg [31:0] _T_574_re; // @[Reg.scala 15:16]
  reg [31:0] _T_574_im; // @[Reg.scala 15:16]
  reg [31:0] _T_575_re; // @[Reg.scala 15:16]
  reg [31:0] _T_575_im; // @[Reg.scala 15:16]
  reg [31:0] _T_576_re; // @[Reg.scala 15:16]
  reg [31:0] _T_576_im; // @[Reg.scala 15:16]
  reg [31:0] _T_577_re; // @[Reg.scala 15:16]
  reg [31:0] _T_577_im; // @[Reg.scala 15:16]
  reg [31:0] _T_578_re; // @[Reg.scala 15:16]
  reg [31:0] _T_578_im; // @[Reg.scala 15:16]
  reg [31:0] _T_579_re; // @[Reg.scala 15:16]
  reg [31:0] _T_579_im; // @[Reg.scala 15:16]
  reg [31:0] _T_580_re; // @[Reg.scala 15:16]
  reg [31:0] _T_580_im; // @[Reg.scala 15:16]
  reg [31:0] _T_581_re; // @[Reg.scala 15:16]
  reg [31:0] _T_581_im; // @[Reg.scala 15:16]
  reg [31:0] _T_582_re; // @[Reg.scala 15:16]
  reg [31:0] _T_582_im; // @[Reg.scala 15:16]
  reg [31:0] _T_583_re; // @[Reg.scala 15:16]
  reg [31:0] _T_583_im; // @[Reg.scala 15:16]
  reg [31:0] _T_584_re; // @[Reg.scala 15:16]
  reg [31:0] _T_584_im; // @[Reg.scala 15:16]
  reg [31:0] _T_585_re; // @[Reg.scala 15:16]
  reg [31:0] _T_585_im; // @[Reg.scala 15:16]
  reg [31:0] _T_586_re; // @[Reg.scala 15:16]
  reg [31:0] _T_586_im; // @[Reg.scala 15:16]
  reg [31:0] _T_587_re; // @[Reg.scala 15:16]
  reg [31:0] _T_587_im; // @[Reg.scala 15:16]
  reg [31:0] _T_588_re; // @[Reg.scala 15:16]
  reg [31:0] _T_588_im; // @[Reg.scala 15:16]
  reg [31:0] _T_589_re; // @[Reg.scala 15:16]
  reg [31:0] _T_589_im; // @[Reg.scala 15:16]
  reg [31:0] _T_590_re; // @[Reg.scala 15:16]
  reg [31:0] _T_590_im; // @[Reg.scala 15:16]
  reg [31:0] _T_591_re; // @[Reg.scala 15:16]
  reg [31:0] _T_591_im; // @[Reg.scala 15:16]
  reg [31:0] _T_592_re; // @[Reg.scala 15:16]
  reg [31:0] _T_592_im; // @[Reg.scala 15:16]
  reg [31:0] _T_593_re; // @[Reg.scala 15:16]
  reg [31:0] _T_593_im; // @[Reg.scala 15:16]
  reg [31:0] _T_594_re; // @[Reg.scala 15:16]
  reg [31:0] _T_594_im; // @[Reg.scala 15:16]
  reg [31:0] _T_595_re; // @[Reg.scala 15:16]
  reg [31:0] _T_595_im; // @[Reg.scala 15:16]
  reg [31:0] _T_596_re; // @[Reg.scala 15:16]
  reg [31:0] _T_596_im; // @[Reg.scala 15:16]
  reg [31:0] _T_597_re; // @[Reg.scala 15:16]
  reg [31:0] _T_597_im; // @[Reg.scala 15:16]
  reg [31:0] _T_598_re; // @[Reg.scala 15:16]
  reg [31:0] _T_598_im; // @[Reg.scala 15:16]
  reg [31:0] _T_599_re; // @[Reg.scala 15:16]
  reg [31:0] _T_599_im; // @[Reg.scala 15:16]
  reg [31:0] _T_600_re; // @[Reg.scala 15:16]
  reg [31:0] _T_600_im; // @[Reg.scala 15:16]
  reg [31:0] _T_601_re; // @[Reg.scala 15:16]
  reg [31:0] _T_601_im; // @[Reg.scala 15:16]
  reg [31:0] _T_602_re; // @[Reg.scala 15:16]
  reg [31:0] _T_602_im; // @[Reg.scala 15:16]
  reg [31:0] _T_603_re; // @[Reg.scala 15:16]
  reg [31:0] _T_603_im; // @[Reg.scala 15:16]
  reg [31:0] _T_604_re; // @[Reg.scala 15:16]
  reg [31:0] _T_604_im; // @[Reg.scala 15:16]
  reg [31:0] _T_605_re; // @[Reg.scala 15:16]
  reg [31:0] _T_605_im; // @[Reg.scala 15:16]
  reg [31:0] _T_606_re; // @[Reg.scala 15:16]
  reg [31:0] _T_606_im; // @[Reg.scala 15:16]
  reg [31:0] _T_607_re; // @[Reg.scala 15:16]
  reg [31:0] _T_607_im; // @[Reg.scala 15:16]
  reg [31:0] _T_608_re; // @[Reg.scala 15:16]
  reg [31:0] _T_608_im; // @[Reg.scala 15:16]
  reg [31:0] _T_609_re; // @[Reg.scala 15:16]
  reg [31:0] _T_609_im; // @[Reg.scala 15:16]
  reg [31:0] _T_610_re; // @[Reg.scala 15:16]
  reg [31:0] _T_610_im; // @[Reg.scala 15:16]
  reg [31:0] _T_611_re; // @[Reg.scala 15:16]
  reg [31:0] _T_611_im; // @[Reg.scala 15:16]
  reg [31:0] _T_612_re; // @[Reg.scala 15:16]
  reg [31:0] _T_612_im; // @[Reg.scala 15:16]
  reg [31:0] _T_613_re; // @[Reg.scala 15:16]
  reg [31:0] _T_613_im; // @[Reg.scala 15:16]
  reg [31:0] _T_614_re; // @[Reg.scala 15:16]
  reg [31:0] _T_614_im; // @[Reg.scala 15:16]
  reg [31:0] _T_615_re; // @[Reg.scala 15:16]
  reg [31:0] _T_615_im; // @[Reg.scala 15:16]
  reg [31:0] _T_616_re; // @[Reg.scala 15:16]
  reg [31:0] _T_616_im; // @[Reg.scala 15:16]
  reg [31:0] _T_617_re; // @[Reg.scala 15:16]
  reg [31:0] _T_617_im; // @[Reg.scala 15:16]
  reg [31:0] _T_618_re; // @[Reg.scala 15:16]
  reg [31:0] _T_618_im; // @[Reg.scala 15:16]
  reg [31:0] _T_619_re; // @[Reg.scala 15:16]
  reg [31:0] _T_619_im; // @[Reg.scala 15:16]
  reg [31:0] _T_620_re; // @[Reg.scala 15:16]
  reg [31:0] _T_620_im; // @[Reg.scala 15:16]
  reg [31:0] _T_621_re; // @[Reg.scala 15:16]
  reg [31:0] _T_621_im; // @[Reg.scala 15:16]
  reg [31:0] _T_622_re; // @[Reg.scala 15:16]
  reg [31:0] _T_622_im; // @[Reg.scala 15:16]
  reg [31:0] _T_623_re; // @[Reg.scala 15:16]
  reg [31:0] _T_623_im; // @[Reg.scala 15:16]
  reg [31:0] _T_624_re; // @[Reg.scala 15:16]
  reg [31:0] _T_624_im; // @[Reg.scala 15:16]
  reg [31:0] _T_625_re; // @[Reg.scala 15:16]
  reg [31:0] _T_625_im; // @[Reg.scala 15:16]
  reg [31:0] _T_626_re; // @[Reg.scala 15:16]
  reg [31:0] _T_626_im; // @[Reg.scala 15:16]
  reg [31:0] _T_627_re; // @[Reg.scala 15:16]
  reg [31:0] _T_627_im; // @[Reg.scala 15:16]
  reg [31:0] _T_628_re; // @[Reg.scala 15:16]
  reg [31:0] _T_628_im; // @[Reg.scala 15:16]
  reg [31:0] _T_629_re; // @[Reg.scala 15:16]
  reg [31:0] _T_629_im; // @[Reg.scala 15:16]
  reg [31:0] _T_630_re; // @[Reg.scala 15:16]
  reg [31:0] _T_630_im; // @[Reg.scala 15:16]
  reg [31:0] _T_631_re; // @[Reg.scala 15:16]
  reg [31:0] _T_631_im; // @[Reg.scala 15:16]
  reg [31:0] _T_632_re; // @[Reg.scala 15:16]
  reg [31:0] _T_632_im; // @[Reg.scala 15:16]
  reg [31:0] _T_633_re; // @[Reg.scala 15:16]
  reg [31:0] _T_633_im; // @[Reg.scala 15:16]
  reg [31:0] _T_634_re; // @[Reg.scala 15:16]
  reg [31:0] _T_634_im; // @[Reg.scala 15:16]
  reg [31:0] _T_635_re; // @[Reg.scala 15:16]
  reg [31:0] _T_635_im; // @[Reg.scala 15:16]
  reg [31:0] _T_636_re; // @[Reg.scala 15:16]
  reg [31:0] _T_636_im; // @[Reg.scala 15:16]
  reg [31:0] _T_637_re; // @[Reg.scala 15:16]
  reg [31:0] _T_637_im; // @[Reg.scala 15:16]
  reg [31:0] _T_638_re; // @[Reg.scala 15:16]
  reg [31:0] _T_638_im; // @[Reg.scala 15:16]
  reg [31:0] _T_639_re; // @[Reg.scala 15:16]
  reg [31:0] _T_639_im; // @[Reg.scala 15:16]
  reg [31:0] _T_640_re; // @[Reg.scala 15:16]
  reg [31:0] _T_640_im; // @[Reg.scala 15:16]
  reg [31:0] _T_641_re; // @[Reg.scala 15:16]
  reg [31:0] _T_641_im; // @[Reg.scala 15:16]
  reg [31:0] _T_642_re; // @[Reg.scala 15:16]
  reg [31:0] _T_642_im; // @[Reg.scala 15:16]
  reg [31:0] _T_643_re; // @[Reg.scala 15:16]
  reg [31:0] _T_643_im; // @[Reg.scala 15:16]
  reg [31:0] _T_644_re; // @[Reg.scala 15:16]
  reg [31:0] _T_644_im; // @[Reg.scala 15:16]
  reg [31:0] _T_645_re; // @[Reg.scala 15:16]
  reg [31:0] _T_645_im; // @[Reg.scala 15:16]
  reg [31:0] _T_646_re; // @[Reg.scala 15:16]
  reg [31:0] _T_646_im; // @[Reg.scala 15:16]
  reg [31:0] _T_647_re; // @[Reg.scala 15:16]
  reg [31:0] _T_647_im; // @[Reg.scala 15:16]
  reg [31:0] _T_648_re; // @[Reg.scala 15:16]
  reg [31:0] _T_648_im; // @[Reg.scala 15:16]
  reg [31:0] _T_649_re; // @[Reg.scala 15:16]
  reg [31:0] _T_649_im; // @[Reg.scala 15:16]
  reg [31:0] _T_650_re; // @[Reg.scala 15:16]
  reg [31:0] _T_650_im; // @[Reg.scala 15:16]
  reg [31:0] _T_651_re; // @[Reg.scala 15:16]
  reg [31:0] _T_651_im; // @[Reg.scala 15:16]
  reg [31:0] _T_652_re; // @[Reg.scala 15:16]
  reg [31:0] _T_652_im; // @[Reg.scala 15:16]
  reg [31:0] _T_653_re; // @[Reg.scala 15:16]
  reg [31:0] _T_653_im; // @[Reg.scala 15:16]
  reg [31:0] _T_654_re; // @[Reg.scala 15:16]
  reg [31:0] _T_654_im; // @[Reg.scala 15:16]
  reg [31:0] _T_655_re; // @[Reg.scala 15:16]
  reg [31:0] _T_655_im; // @[Reg.scala 15:16]
  reg [31:0] _T_656_re; // @[Reg.scala 15:16]
  reg [31:0] _T_656_im; // @[Reg.scala 15:16]
  reg [31:0] _T_657_re; // @[Reg.scala 15:16]
  reg [31:0] _T_657_im; // @[Reg.scala 15:16]
  reg [31:0] _T_658_re; // @[Reg.scala 15:16]
  reg [31:0] _T_658_im; // @[Reg.scala 15:16]
  reg [31:0] _T_659_re; // @[Reg.scala 15:16]
  reg [31:0] _T_659_im; // @[Reg.scala 15:16]
  reg [31:0] _T_660_re; // @[Reg.scala 15:16]
  reg [31:0] _T_660_im; // @[Reg.scala 15:16]
  reg [31:0] _T_661_re; // @[Reg.scala 15:16]
  reg [31:0] _T_661_im; // @[Reg.scala 15:16]
  reg [31:0] _T_662_re; // @[Reg.scala 15:16]
  reg [31:0] _T_662_im; // @[Reg.scala 15:16]
  reg [31:0] _T_663_re; // @[Reg.scala 15:16]
  reg [31:0] _T_663_im; // @[Reg.scala 15:16]
  reg [31:0] _T_664_re; // @[Reg.scala 15:16]
  reg [31:0] _T_664_im; // @[Reg.scala 15:16]
  reg [31:0] _T_665_re; // @[Reg.scala 15:16]
  reg [31:0] _T_665_im; // @[Reg.scala 15:16]
  reg [31:0] _T_666_re; // @[Reg.scala 15:16]
  reg [31:0] _T_666_im; // @[Reg.scala 15:16]
  reg [31:0] _T_667_re; // @[Reg.scala 15:16]
  reg [31:0] _T_667_im; // @[Reg.scala 15:16]
  reg [31:0] _T_668_re; // @[Reg.scala 15:16]
  reg [31:0] _T_668_im; // @[Reg.scala 15:16]
  reg [31:0] _T_669_re; // @[Reg.scala 15:16]
  reg [31:0] _T_669_im; // @[Reg.scala 15:16]
  reg [31:0] _T_670_re; // @[Reg.scala 15:16]
  reg [31:0] _T_670_im; // @[Reg.scala 15:16]
  reg [31:0] _T_672_re; // @[Reg.scala 15:16]
  reg [31:0] _T_672_im; // @[Reg.scala 15:16]
  reg [31:0] _T_673_re; // @[Reg.scala 15:16]
  reg [31:0] _T_673_im; // @[Reg.scala 15:16]
  reg [31:0] _T_674_re; // @[Reg.scala 15:16]
  reg [31:0] _T_674_im; // @[Reg.scala 15:16]
  reg [31:0] _T_675_re; // @[Reg.scala 15:16]
  reg [31:0] _T_675_im; // @[Reg.scala 15:16]
  reg [31:0] _T_676_re; // @[Reg.scala 15:16]
  reg [31:0] _T_676_im; // @[Reg.scala 15:16]
  reg [31:0] _T_677_re; // @[Reg.scala 15:16]
  reg [31:0] _T_677_im; // @[Reg.scala 15:16]
  reg [31:0] _T_678_re; // @[Reg.scala 15:16]
  reg [31:0] _T_678_im; // @[Reg.scala 15:16]
  reg [31:0] _T_679_re; // @[Reg.scala 15:16]
  reg [31:0] _T_679_im; // @[Reg.scala 15:16]
  reg [31:0] _T_680_re; // @[Reg.scala 15:16]
  reg [31:0] _T_680_im; // @[Reg.scala 15:16]
  reg [31:0] _T_681_re; // @[Reg.scala 15:16]
  reg [31:0] _T_681_im; // @[Reg.scala 15:16]
  reg [31:0] _T_682_re; // @[Reg.scala 15:16]
  reg [31:0] _T_682_im; // @[Reg.scala 15:16]
  reg [31:0] _T_683_re; // @[Reg.scala 15:16]
  reg [31:0] _T_683_im; // @[Reg.scala 15:16]
  reg [31:0] _T_684_re; // @[Reg.scala 15:16]
  reg [31:0] _T_684_im; // @[Reg.scala 15:16]
  reg [31:0] _T_685_re; // @[Reg.scala 15:16]
  reg [31:0] _T_685_im; // @[Reg.scala 15:16]
  reg [31:0] _T_686_re; // @[Reg.scala 15:16]
  reg [31:0] _T_686_im; // @[Reg.scala 15:16]
  reg [31:0] _T_687_re; // @[Reg.scala 15:16]
  reg [31:0] _T_687_im; // @[Reg.scala 15:16]
  reg [31:0] _T_688_re; // @[Reg.scala 15:16]
  reg [31:0] _T_688_im; // @[Reg.scala 15:16]
  reg [31:0] _T_689_re; // @[Reg.scala 15:16]
  reg [31:0] _T_689_im; // @[Reg.scala 15:16]
  reg [31:0] _T_690_re; // @[Reg.scala 15:16]
  reg [31:0] _T_690_im; // @[Reg.scala 15:16]
  reg [31:0] _T_691_re; // @[Reg.scala 15:16]
  reg [31:0] _T_691_im; // @[Reg.scala 15:16]
  reg [31:0] _T_692_re; // @[Reg.scala 15:16]
  reg [31:0] _T_692_im; // @[Reg.scala 15:16]
  reg [31:0] _T_693_re; // @[Reg.scala 15:16]
  reg [31:0] _T_693_im; // @[Reg.scala 15:16]
  reg [31:0] _T_694_re; // @[Reg.scala 15:16]
  reg [31:0] _T_694_im; // @[Reg.scala 15:16]
  reg [31:0] _T_695_re; // @[Reg.scala 15:16]
  reg [31:0] _T_695_im; // @[Reg.scala 15:16]
  reg [31:0] _T_696_re; // @[Reg.scala 15:16]
  reg [31:0] _T_696_im; // @[Reg.scala 15:16]
  reg [31:0] _T_697_re; // @[Reg.scala 15:16]
  reg [31:0] _T_697_im; // @[Reg.scala 15:16]
  reg [31:0] _T_698_re; // @[Reg.scala 15:16]
  reg [31:0] _T_698_im; // @[Reg.scala 15:16]
  reg [31:0] _T_699_re; // @[Reg.scala 15:16]
  reg [31:0] _T_699_im; // @[Reg.scala 15:16]
  reg [31:0] _T_700_re; // @[Reg.scala 15:16]
  reg [31:0] _T_700_im; // @[Reg.scala 15:16]
  reg [31:0] _T_701_re; // @[Reg.scala 15:16]
  reg [31:0] _T_701_im; // @[Reg.scala 15:16]
  reg [31:0] _T_702_re; // @[Reg.scala 15:16]
  reg [31:0] _T_702_im; // @[Reg.scala 15:16]
  reg [31:0] _T_703_re; // @[Reg.scala 15:16]
  reg [31:0] _T_703_im; // @[Reg.scala 15:16]
  reg [31:0] _T_704_re; // @[Reg.scala 15:16]
  reg [31:0] _T_704_im; // @[Reg.scala 15:16]
  reg [31:0] _T_705_re; // @[Reg.scala 15:16]
  reg [31:0] _T_705_im; // @[Reg.scala 15:16]
  reg [31:0] _T_706_re; // @[Reg.scala 15:16]
  reg [31:0] _T_706_im; // @[Reg.scala 15:16]
  reg [31:0] _T_707_re; // @[Reg.scala 15:16]
  reg [31:0] _T_707_im; // @[Reg.scala 15:16]
  reg [31:0] _T_708_re; // @[Reg.scala 15:16]
  reg [31:0] _T_708_im; // @[Reg.scala 15:16]
  reg [31:0] _T_709_re; // @[Reg.scala 15:16]
  reg [31:0] _T_709_im; // @[Reg.scala 15:16]
  reg [31:0] _T_710_re; // @[Reg.scala 15:16]
  reg [31:0] _T_710_im; // @[Reg.scala 15:16]
  reg [31:0] _T_711_re; // @[Reg.scala 15:16]
  reg [31:0] _T_711_im; // @[Reg.scala 15:16]
  reg [31:0] _T_712_re; // @[Reg.scala 15:16]
  reg [31:0] _T_712_im; // @[Reg.scala 15:16]
  reg [31:0] _T_713_re; // @[Reg.scala 15:16]
  reg [31:0] _T_713_im; // @[Reg.scala 15:16]
  reg [31:0] _T_714_re; // @[Reg.scala 15:16]
  reg [31:0] _T_714_im; // @[Reg.scala 15:16]
  reg [31:0] _T_715_re; // @[Reg.scala 15:16]
  reg [31:0] _T_715_im; // @[Reg.scala 15:16]
  reg [31:0] _T_716_re; // @[Reg.scala 15:16]
  reg [31:0] _T_716_im; // @[Reg.scala 15:16]
  reg [31:0] _T_717_re; // @[Reg.scala 15:16]
  reg [31:0] _T_717_im; // @[Reg.scala 15:16]
  reg [31:0] _T_718_re; // @[Reg.scala 15:16]
  reg [31:0] _T_718_im; // @[Reg.scala 15:16]
  reg [31:0] _T_719_re; // @[Reg.scala 15:16]
  reg [31:0] _T_719_im; // @[Reg.scala 15:16]
  reg [31:0] _T_720_re; // @[Reg.scala 15:16]
  reg [31:0] _T_720_im; // @[Reg.scala 15:16]
  reg [31:0] _T_721_re; // @[Reg.scala 15:16]
  reg [31:0] _T_721_im; // @[Reg.scala 15:16]
  reg [31:0] _T_722_re; // @[Reg.scala 15:16]
  reg [31:0] _T_722_im; // @[Reg.scala 15:16]
  reg [31:0] _T_723_re; // @[Reg.scala 15:16]
  reg [31:0] _T_723_im; // @[Reg.scala 15:16]
  reg [31:0] _T_724_re; // @[Reg.scala 15:16]
  reg [31:0] _T_724_im; // @[Reg.scala 15:16]
  reg [31:0] _T_725_re; // @[Reg.scala 15:16]
  reg [31:0] _T_725_im; // @[Reg.scala 15:16]
  reg [31:0] _T_726_re; // @[Reg.scala 15:16]
  reg [31:0] _T_726_im; // @[Reg.scala 15:16]
  reg [31:0] _T_727_re; // @[Reg.scala 15:16]
  reg [31:0] _T_727_im; // @[Reg.scala 15:16]
  reg [31:0] _T_728_re; // @[Reg.scala 15:16]
  reg [31:0] _T_728_im; // @[Reg.scala 15:16]
  reg [31:0] _T_729_re; // @[Reg.scala 15:16]
  reg [31:0] _T_729_im; // @[Reg.scala 15:16]
  reg [31:0] _T_730_re; // @[Reg.scala 15:16]
  reg [31:0] _T_730_im; // @[Reg.scala 15:16]
  reg [31:0] _T_731_re; // @[Reg.scala 15:16]
  reg [31:0] _T_731_im; // @[Reg.scala 15:16]
  reg [31:0] _T_732_re; // @[Reg.scala 15:16]
  reg [31:0] _T_732_im; // @[Reg.scala 15:16]
  reg [31:0] _T_733_re; // @[Reg.scala 15:16]
  reg [31:0] _T_733_im; // @[Reg.scala 15:16]
  reg [31:0] _T_734_re; // @[Reg.scala 15:16]
  reg [31:0] _T_734_im; // @[Reg.scala 15:16]
  reg [31:0] _T_735_re; // @[Reg.scala 15:16]
  reg [31:0] _T_735_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_2690 = 6'h1 == cnt[5:0] ? $signed(32'shffb1) : $signed(32'sh10000); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2691 = 6'h2 == cnt[5:0] ? $signed(32'shfec4) : $signed(_GEN_2690); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2692 = 6'h3 == cnt[5:0] ? $signed(32'shfd3b) : $signed(_GEN_2691); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2693 = 6'h4 == cnt[5:0] ? $signed(32'shfb15) : $signed(_GEN_2692); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2694 = 6'h5 == cnt[5:0] ? $signed(32'shf854) : $signed(_GEN_2693); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2695 = 6'h6 == cnt[5:0] ? $signed(32'shf4fa) : $signed(_GEN_2694); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2696 = 6'h7 == cnt[5:0] ? $signed(32'shf109) : $signed(_GEN_2695); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2697 = 6'h8 == cnt[5:0] ? $signed(32'shec83) : $signed(_GEN_2696); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2698 = 6'h9 == cnt[5:0] ? $signed(32'she76c) : $signed(_GEN_2697); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2699 = 6'ha == cnt[5:0] ? $signed(32'she1c6) : $signed(_GEN_2698); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2700 = 6'hb == cnt[5:0] ? $signed(32'shdb94) : $signed(_GEN_2699); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2701 = 6'hc == cnt[5:0] ? $signed(32'shd4db) : $signed(_GEN_2700); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2702 = 6'hd == cnt[5:0] ? $signed(32'shcd9f) : $signed(_GEN_2701); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2703 = 6'he == cnt[5:0] ? $signed(32'shc5e4) : $signed(_GEN_2702); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2704 = 6'hf == cnt[5:0] ? $signed(32'shbdaf) : $signed(_GEN_2703); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2705 = 6'h10 == cnt[5:0] ? $signed(32'shb505) : $signed(_GEN_2704); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2706 = 6'h11 == cnt[5:0] ? $signed(32'shabeb) : $signed(_GEN_2705); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2707 = 6'h12 == cnt[5:0] ? $signed(32'sha268) : $signed(_GEN_2706); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2708 = 6'h13 == cnt[5:0] ? $signed(32'sh9880) : $signed(_GEN_2707); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2709 = 6'h14 == cnt[5:0] ? $signed(32'sh8e3a) : $signed(_GEN_2708); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2710 = 6'h15 == cnt[5:0] ? $signed(32'sh839c) : $signed(_GEN_2709); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2711 = 6'h16 == cnt[5:0] ? $signed(32'sh78ad) : $signed(_GEN_2710); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2712 = 6'h17 == cnt[5:0] ? $signed(32'sh6d74) : $signed(_GEN_2711); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2713 = 6'h18 == cnt[5:0] ? $signed(32'sh61f8) : $signed(_GEN_2712); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2714 = 6'h19 == cnt[5:0] ? $signed(32'sh563e) : $signed(_GEN_2713); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2715 = 6'h1a == cnt[5:0] ? $signed(32'sh4a50) : $signed(_GEN_2714); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2716 = 6'h1b == cnt[5:0] ? $signed(32'sh3e34) : $signed(_GEN_2715); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2717 = 6'h1c == cnt[5:0] ? $signed(32'sh31f1) : $signed(_GEN_2716); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2718 = 6'h1d == cnt[5:0] ? $signed(32'sh2590) : $signed(_GEN_2717); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2719 = 6'h1e == cnt[5:0] ? $signed(32'sh1918) : $signed(_GEN_2718); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2720 = 6'h1f == cnt[5:0] ? $signed(32'shc90) : $signed(_GEN_2719); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2721 = 6'h20 == cnt[5:0] ? $signed(32'sh0) : $signed(_GEN_2720); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2722 = 6'h21 == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_2721); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2723 = 6'h22 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_2722); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2724 = 6'h23 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_2723); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2725 = 6'h24 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_2724); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2726 = 6'h25 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_2725); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2727 = 6'h26 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_2726); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2728 = 6'h27 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_2727); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2729 = 6'h28 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_2728); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2730 = 6'h29 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_2729); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2731 = 6'h2a == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_2730); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2732 = 6'h2b == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_2731); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2733 = 6'h2c == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2732); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2734 = 6'h2d == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_2733); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2735 = 6'h2e == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_2734); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2736 = 6'h2f == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_2735); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2737 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2736); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2738 = 6'h31 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2737); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2739 = 6'h32 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2738); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2740 = 6'h33 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2739); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2741 = 6'h34 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2740); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2742 = 6'h35 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2741); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2743 = 6'h36 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2742); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2744 = 6'h37 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2743); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2745 = 6'h38 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2744); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2746 = 6'h39 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2745); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2747 = 6'h3a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2746); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2748 = 6'h3b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2747); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2749 = 6'h3c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2748); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2750 = 6'h3d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2749); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2751 = 6'h3e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2750); // @[FFT.scala 51:18]
  wire [31:0] _GEN_2882 = 6'h1 == cnt[5:0] ? $signed(-32'shc90) : $signed(32'sh0); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2883 = 6'h2 == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_2882); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2884 = 6'h3 == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_2883); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2885 = 6'h4 == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_2884); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2886 = 6'h5 == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_2885); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2887 = 6'h6 == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_2886); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2888 = 6'h7 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_2887); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2889 = 6'h8 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_2888); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2890 = 6'h9 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_2889); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2891 = 6'ha == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_2890); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2892 = 6'hb == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_2891); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2893 = 6'hc == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2892); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2894 = 6'hd == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_2893); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2895 = 6'he == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_2894); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2896 = 6'hf == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_2895); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2897 = 6'h10 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2896); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2898 = 6'h11 == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2897); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2899 = 6'h12 == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2898); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2900 = 6'h13 == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2899); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2901 = 6'h14 == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2900); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2902 = 6'h15 == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2901); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2903 = 6'h16 == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2902); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2904 = 6'h17 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2903); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2905 = 6'h18 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2904); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2906 = 6'h19 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2905); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2907 = 6'h1a == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2906); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2908 = 6'h1b == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2907); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2909 = 6'h1c == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2908); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2910 = 6'h1d == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2909); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2911 = 6'h1e == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2910); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2912 = 6'h1f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2911); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2913 = 6'h20 == cnt[5:0] ? $signed(-32'sh10000) : $signed(_GEN_2912); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2914 = 6'h21 == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2913); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2915 = 6'h22 == cnt[5:0] ? $signed(-32'shfec4) : $signed(_GEN_2914); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2916 = 6'h23 == cnt[5:0] ? $signed(-32'shfd3b) : $signed(_GEN_2915); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2917 = 6'h24 == cnt[5:0] ? $signed(-32'shfb15) : $signed(_GEN_2916); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2918 = 6'h25 == cnt[5:0] ? $signed(-32'shf854) : $signed(_GEN_2917); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2919 = 6'h26 == cnt[5:0] ? $signed(-32'shf4fa) : $signed(_GEN_2918); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2920 = 6'h27 == cnt[5:0] ? $signed(-32'shf109) : $signed(_GEN_2919); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2921 = 6'h28 == cnt[5:0] ? $signed(-32'shec83) : $signed(_GEN_2920); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2922 = 6'h29 == cnt[5:0] ? $signed(-32'she76c) : $signed(_GEN_2921); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2923 = 6'h2a == cnt[5:0] ? $signed(-32'she1c6) : $signed(_GEN_2922); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2924 = 6'h2b == cnt[5:0] ? $signed(-32'shdb94) : $signed(_GEN_2923); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2925 = 6'h2c == cnt[5:0] ? $signed(-32'shd4db) : $signed(_GEN_2924); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2926 = 6'h2d == cnt[5:0] ? $signed(-32'shcd9f) : $signed(_GEN_2925); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2927 = 6'h2e == cnt[5:0] ? $signed(-32'shc5e4) : $signed(_GEN_2926); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2928 = 6'h2f == cnt[5:0] ? $signed(-32'shbdaf) : $signed(_GEN_2927); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2929 = 6'h30 == cnt[5:0] ? $signed(-32'shb505) : $signed(_GEN_2928); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2930 = 6'h31 == cnt[5:0] ? $signed(-32'shabeb) : $signed(_GEN_2929); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2931 = 6'h32 == cnt[5:0] ? $signed(-32'sha268) : $signed(_GEN_2930); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2932 = 6'h33 == cnt[5:0] ? $signed(-32'sh9880) : $signed(_GEN_2931); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2933 = 6'h34 == cnt[5:0] ? $signed(-32'sh8e3a) : $signed(_GEN_2932); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2934 = 6'h35 == cnt[5:0] ? $signed(-32'sh839c) : $signed(_GEN_2933); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2935 = 6'h36 == cnt[5:0] ? $signed(-32'sh78ad) : $signed(_GEN_2934); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2936 = 6'h37 == cnt[5:0] ? $signed(-32'sh6d74) : $signed(_GEN_2935); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2937 = 6'h38 == cnt[5:0] ? $signed(-32'sh61f8) : $signed(_GEN_2936); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2938 = 6'h39 == cnt[5:0] ? $signed(-32'sh563e) : $signed(_GEN_2937); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2939 = 6'h3a == cnt[5:0] ? $signed(-32'sh4a50) : $signed(_GEN_2938); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2940 = 6'h3b == cnt[5:0] ? $signed(-32'sh3e34) : $signed(_GEN_2939); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2941 = 6'h3c == cnt[5:0] ? $signed(-32'sh31f1) : $signed(_GEN_2940); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2942 = 6'h3d == cnt[5:0] ? $signed(-32'sh2590) : $signed(_GEN_2941); // @[FFT.scala 52:18]
  wire [31:0] _GEN_2943 = 6'h3e == cnt[5:0] ? $signed(-32'sh1918) : $signed(_GEN_2942); // @[FFT.scala 52:18]
  reg [31:0] _T_744_re; // @[Reg.scala 15:16]
  reg [31:0] _T_744_im; // @[Reg.scala 15:16]
  reg [31:0] _T_745_re; // @[Reg.scala 15:16]
  reg [31:0] _T_745_im; // @[Reg.scala 15:16]
  reg [31:0] _T_746_re; // @[Reg.scala 15:16]
  reg [31:0] _T_746_im; // @[Reg.scala 15:16]
  reg [31:0] _T_747_re; // @[Reg.scala 15:16]
  reg [31:0] _T_747_im; // @[Reg.scala 15:16]
  reg [31:0] _T_748_re; // @[Reg.scala 15:16]
  reg [31:0] _T_748_im; // @[Reg.scala 15:16]
  reg [31:0] _T_749_re; // @[Reg.scala 15:16]
  reg [31:0] _T_749_im; // @[Reg.scala 15:16]
  reg [31:0] _T_750_re; // @[Reg.scala 15:16]
  reg [31:0] _T_750_im; // @[Reg.scala 15:16]
  reg [31:0] _T_751_re; // @[Reg.scala 15:16]
  reg [31:0] _T_751_im; // @[Reg.scala 15:16]
  reg [31:0] _T_752_re; // @[Reg.scala 15:16]
  reg [31:0] _T_752_im; // @[Reg.scala 15:16]
  reg [31:0] _T_753_re; // @[Reg.scala 15:16]
  reg [31:0] _T_753_im; // @[Reg.scala 15:16]
  reg [31:0] _T_754_re; // @[Reg.scala 15:16]
  reg [31:0] _T_754_im; // @[Reg.scala 15:16]
  reg [31:0] _T_755_re; // @[Reg.scala 15:16]
  reg [31:0] _T_755_im; // @[Reg.scala 15:16]
  reg [31:0] _T_756_re; // @[Reg.scala 15:16]
  reg [31:0] _T_756_im; // @[Reg.scala 15:16]
  reg [31:0] _T_757_re; // @[Reg.scala 15:16]
  reg [31:0] _T_757_im; // @[Reg.scala 15:16]
  reg [31:0] _T_758_re; // @[Reg.scala 15:16]
  reg [31:0] _T_758_im; // @[Reg.scala 15:16]
  reg [31:0] _T_759_re; // @[Reg.scala 15:16]
  reg [31:0] _T_759_im; // @[Reg.scala 15:16]
  reg [31:0] _T_760_re; // @[Reg.scala 15:16]
  reg [31:0] _T_760_im; // @[Reg.scala 15:16]
  reg [31:0] _T_761_re; // @[Reg.scala 15:16]
  reg [31:0] _T_761_im; // @[Reg.scala 15:16]
  reg [31:0] _T_762_re; // @[Reg.scala 15:16]
  reg [31:0] _T_762_im; // @[Reg.scala 15:16]
  reg [31:0] _T_763_re; // @[Reg.scala 15:16]
  reg [31:0] _T_763_im; // @[Reg.scala 15:16]
  reg [31:0] _T_764_re; // @[Reg.scala 15:16]
  reg [31:0] _T_764_im; // @[Reg.scala 15:16]
  reg [31:0] _T_765_re; // @[Reg.scala 15:16]
  reg [31:0] _T_765_im; // @[Reg.scala 15:16]
  reg [31:0] _T_766_re; // @[Reg.scala 15:16]
  reg [31:0] _T_766_im; // @[Reg.scala 15:16]
  reg [31:0] _T_767_re; // @[Reg.scala 15:16]
  reg [31:0] _T_767_im; // @[Reg.scala 15:16]
  reg [31:0] _T_768_re; // @[Reg.scala 15:16]
  reg [31:0] _T_768_im; // @[Reg.scala 15:16]
  reg [31:0] _T_769_re; // @[Reg.scala 15:16]
  reg [31:0] _T_769_im; // @[Reg.scala 15:16]
  reg [31:0] _T_770_re; // @[Reg.scala 15:16]
  reg [31:0] _T_770_im; // @[Reg.scala 15:16]
  reg [31:0] _T_771_re; // @[Reg.scala 15:16]
  reg [31:0] _T_771_im; // @[Reg.scala 15:16]
  reg [31:0] _T_772_re; // @[Reg.scala 15:16]
  reg [31:0] _T_772_im; // @[Reg.scala 15:16]
  reg [31:0] _T_773_re; // @[Reg.scala 15:16]
  reg [31:0] _T_773_im; // @[Reg.scala 15:16]
  reg [31:0] _T_774_re; // @[Reg.scala 15:16]
  reg [31:0] _T_774_im; // @[Reg.scala 15:16]
  reg [31:0] _T_775_re; // @[Reg.scala 15:16]
  reg [31:0] _T_775_im; // @[Reg.scala 15:16]
  reg [31:0] _T_776_re; // @[Reg.scala 15:16]
  reg [31:0] _T_776_im; // @[Reg.scala 15:16]
  reg [31:0] _T_777_re; // @[Reg.scala 15:16]
  reg [31:0] _T_777_im; // @[Reg.scala 15:16]
  reg [31:0] _T_778_re; // @[Reg.scala 15:16]
  reg [31:0] _T_778_im; // @[Reg.scala 15:16]
  reg [31:0] _T_779_re; // @[Reg.scala 15:16]
  reg [31:0] _T_779_im; // @[Reg.scala 15:16]
  reg [31:0] _T_780_re; // @[Reg.scala 15:16]
  reg [31:0] _T_780_im; // @[Reg.scala 15:16]
  reg [31:0] _T_781_re; // @[Reg.scala 15:16]
  reg [31:0] _T_781_im; // @[Reg.scala 15:16]
  reg [31:0] _T_782_re; // @[Reg.scala 15:16]
  reg [31:0] _T_782_im; // @[Reg.scala 15:16]
  reg [31:0] _T_783_re; // @[Reg.scala 15:16]
  reg [31:0] _T_783_im; // @[Reg.scala 15:16]
  reg [31:0] _T_784_re; // @[Reg.scala 15:16]
  reg [31:0] _T_784_im; // @[Reg.scala 15:16]
  reg [31:0] _T_785_re; // @[Reg.scala 15:16]
  reg [31:0] _T_785_im; // @[Reg.scala 15:16]
  reg [31:0] _T_786_re; // @[Reg.scala 15:16]
  reg [31:0] _T_786_im; // @[Reg.scala 15:16]
  reg [31:0] _T_787_re; // @[Reg.scala 15:16]
  reg [31:0] _T_787_im; // @[Reg.scala 15:16]
  reg [31:0] _T_788_re; // @[Reg.scala 15:16]
  reg [31:0] _T_788_im; // @[Reg.scala 15:16]
  reg [31:0] _T_789_re; // @[Reg.scala 15:16]
  reg [31:0] _T_789_im; // @[Reg.scala 15:16]
  reg [31:0] _T_790_re; // @[Reg.scala 15:16]
  reg [31:0] _T_790_im; // @[Reg.scala 15:16]
  reg [31:0] _T_791_re; // @[Reg.scala 15:16]
  reg [31:0] _T_791_im; // @[Reg.scala 15:16]
  reg [31:0] _T_792_re; // @[Reg.scala 15:16]
  reg [31:0] _T_792_im; // @[Reg.scala 15:16]
  reg [31:0] _T_793_re; // @[Reg.scala 15:16]
  reg [31:0] _T_793_im; // @[Reg.scala 15:16]
  reg [31:0] _T_794_re; // @[Reg.scala 15:16]
  reg [31:0] _T_794_im; // @[Reg.scala 15:16]
  reg [31:0] _T_795_re; // @[Reg.scala 15:16]
  reg [31:0] _T_795_im; // @[Reg.scala 15:16]
  reg [31:0] _T_796_re; // @[Reg.scala 15:16]
  reg [31:0] _T_796_im; // @[Reg.scala 15:16]
  reg [31:0] _T_797_re; // @[Reg.scala 15:16]
  reg [31:0] _T_797_im; // @[Reg.scala 15:16]
  reg [31:0] _T_798_re; // @[Reg.scala 15:16]
  reg [31:0] _T_798_im; // @[Reg.scala 15:16]
  reg [31:0] _T_799_re; // @[Reg.scala 15:16]
  reg [31:0] _T_799_im; // @[Reg.scala 15:16]
  reg [31:0] _T_800_re; // @[Reg.scala 15:16]
  reg [31:0] _T_800_im; // @[Reg.scala 15:16]
  reg [31:0] _T_801_re; // @[Reg.scala 15:16]
  reg [31:0] _T_801_im; // @[Reg.scala 15:16]
  reg [31:0] _T_802_re; // @[Reg.scala 15:16]
  reg [31:0] _T_802_im; // @[Reg.scala 15:16]
  reg [31:0] _T_803_re; // @[Reg.scala 15:16]
  reg [31:0] _T_803_im; // @[Reg.scala 15:16]
  reg [31:0] _T_804_re; // @[Reg.scala 15:16]
  reg [31:0] _T_804_im; // @[Reg.scala 15:16]
  reg [31:0] _T_805_re; // @[Reg.scala 15:16]
  reg [31:0] _T_805_im; // @[Reg.scala 15:16]
  reg [31:0] _T_806_re; // @[Reg.scala 15:16]
  reg [31:0] _T_806_im; // @[Reg.scala 15:16]
  reg [31:0] _T_807_re; // @[Reg.scala 15:16]
  reg [31:0] _T_807_im; // @[Reg.scala 15:16]
  reg [31:0] _T_809_re; // @[Reg.scala 15:16]
  reg [31:0] _T_809_im; // @[Reg.scala 15:16]
  reg [31:0] _T_810_re; // @[Reg.scala 15:16]
  reg [31:0] _T_810_im; // @[Reg.scala 15:16]
  reg [31:0] _T_811_re; // @[Reg.scala 15:16]
  reg [31:0] _T_811_im; // @[Reg.scala 15:16]
  reg [31:0] _T_812_re; // @[Reg.scala 15:16]
  reg [31:0] _T_812_im; // @[Reg.scala 15:16]
  reg [31:0] _T_813_re; // @[Reg.scala 15:16]
  reg [31:0] _T_813_im; // @[Reg.scala 15:16]
  reg [31:0] _T_814_re; // @[Reg.scala 15:16]
  reg [31:0] _T_814_im; // @[Reg.scala 15:16]
  reg [31:0] _T_815_re; // @[Reg.scala 15:16]
  reg [31:0] _T_815_im; // @[Reg.scala 15:16]
  reg [31:0] _T_816_re; // @[Reg.scala 15:16]
  reg [31:0] _T_816_im; // @[Reg.scala 15:16]
  reg [31:0] _T_817_re; // @[Reg.scala 15:16]
  reg [31:0] _T_817_im; // @[Reg.scala 15:16]
  reg [31:0] _T_818_re; // @[Reg.scala 15:16]
  reg [31:0] _T_818_im; // @[Reg.scala 15:16]
  reg [31:0] _T_819_re; // @[Reg.scala 15:16]
  reg [31:0] _T_819_im; // @[Reg.scala 15:16]
  reg [31:0] _T_820_re; // @[Reg.scala 15:16]
  reg [31:0] _T_820_im; // @[Reg.scala 15:16]
  reg [31:0] _T_821_re; // @[Reg.scala 15:16]
  reg [31:0] _T_821_im; // @[Reg.scala 15:16]
  reg [31:0] _T_822_re; // @[Reg.scala 15:16]
  reg [31:0] _T_822_im; // @[Reg.scala 15:16]
  reg [31:0] _T_823_re; // @[Reg.scala 15:16]
  reg [31:0] _T_823_im; // @[Reg.scala 15:16]
  reg [31:0] _T_824_re; // @[Reg.scala 15:16]
  reg [31:0] _T_824_im; // @[Reg.scala 15:16]
  reg [31:0] _T_825_re; // @[Reg.scala 15:16]
  reg [31:0] _T_825_im; // @[Reg.scala 15:16]
  reg [31:0] _T_826_re; // @[Reg.scala 15:16]
  reg [31:0] _T_826_im; // @[Reg.scala 15:16]
  reg [31:0] _T_827_re; // @[Reg.scala 15:16]
  reg [31:0] _T_827_im; // @[Reg.scala 15:16]
  reg [31:0] _T_828_re; // @[Reg.scala 15:16]
  reg [31:0] _T_828_im; // @[Reg.scala 15:16]
  reg [31:0] _T_829_re; // @[Reg.scala 15:16]
  reg [31:0] _T_829_im; // @[Reg.scala 15:16]
  reg [31:0] _T_830_re; // @[Reg.scala 15:16]
  reg [31:0] _T_830_im; // @[Reg.scala 15:16]
  reg [31:0] _T_831_re; // @[Reg.scala 15:16]
  reg [31:0] _T_831_im; // @[Reg.scala 15:16]
  reg [31:0] _T_832_re; // @[Reg.scala 15:16]
  reg [31:0] _T_832_im; // @[Reg.scala 15:16]
  reg [31:0] _T_833_re; // @[Reg.scala 15:16]
  reg [31:0] _T_833_im; // @[Reg.scala 15:16]
  reg [31:0] _T_834_re; // @[Reg.scala 15:16]
  reg [31:0] _T_834_im; // @[Reg.scala 15:16]
  reg [31:0] _T_835_re; // @[Reg.scala 15:16]
  reg [31:0] _T_835_im; // @[Reg.scala 15:16]
  reg [31:0] _T_836_re; // @[Reg.scala 15:16]
  reg [31:0] _T_836_im; // @[Reg.scala 15:16]
  reg [31:0] _T_837_re; // @[Reg.scala 15:16]
  reg [31:0] _T_837_im; // @[Reg.scala 15:16]
  reg [31:0] _T_838_re; // @[Reg.scala 15:16]
  reg [31:0] _T_838_im; // @[Reg.scala 15:16]
  reg [31:0] _T_839_re; // @[Reg.scala 15:16]
  reg [31:0] _T_839_im; // @[Reg.scala 15:16]
  reg [31:0] _T_840_re; // @[Reg.scala 15:16]
  reg [31:0] _T_840_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3138 = 5'h1 == cnt[4:0] ? $signed(32'shfec4) : $signed(32'sh10000); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3139 = 5'h2 == cnt[4:0] ? $signed(32'shfb15) : $signed(_GEN_3138); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3140 = 5'h3 == cnt[4:0] ? $signed(32'shf4fa) : $signed(_GEN_3139); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3141 = 5'h4 == cnt[4:0] ? $signed(32'shec83) : $signed(_GEN_3140); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3142 = 5'h5 == cnt[4:0] ? $signed(32'she1c6) : $signed(_GEN_3141); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3143 = 5'h6 == cnt[4:0] ? $signed(32'shd4db) : $signed(_GEN_3142); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3144 = 5'h7 == cnt[4:0] ? $signed(32'shc5e4) : $signed(_GEN_3143); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3145 = 5'h8 == cnt[4:0] ? $signed(32'shb505) : $signed(_GEN_3144); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3146 = 5'h9 == cnt[4:0] ? $signed(32'sha268) : $signed(_GEN_3145); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3147 = 5'ha == cnt[4:0] ? $signed(32'sh8e3a) : $signed(_GEN_3146); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3148 = 5'hb == cnt[4:0] ? $signed(32'sh78ad) : $signed(_GEN_3147); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3149 = 5'hc == cnt[4:0] ? $signed(32'sh61f8) : $signed(_GEN_3148); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3150 = 5'hd == cnt[4:0] ? $signed(32'sh4a50) : $signed(_GEN_3149); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3151 = 5'he == cnt[4:0] ? $signed(32'sh31f1) : $signed(_GEN_3150); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3152 = 5'hf == cnt[4:0] ? $signed(32'sh1918) : $signed(_GEN_3151); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3153 = 5'h10 == cnt[4:0] ? $signed(32'sh0) : $signed(_GEN_3152); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3154 = 5'h11 == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_3153); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3155 = 5'h12 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_3154); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3156 = 5'h13 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_3155); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3157 = 5'h14 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_3156); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3158 = 5'h15 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_3157); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3159 = 5'h16 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3158); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3160 = 5'h17 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_3159); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3161 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_3160); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3162 = 5'h19 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_3161); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3163 = 5'h1a == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_3162); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3164 = 5'h1b == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_3163); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3165 = 5'h1c == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_3164); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3166 = 5'h1d == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_3165); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3167 = 5'h1e == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_3166); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3234 = 5'h1 == cnt[4:0] ? $signed(-32'sh1918) : $signed(32'sh0); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3235 = 5'h2 == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_3234); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3236 = 5'h3 == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_3235); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3237 = 5'h4 == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_3236); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3238 = 5'h5 == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_3237); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3239 = 5'h6 == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3238); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3240 = 5'h7 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_3239); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3241 = 5'h8 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_3240); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3242 = 5'h9 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_3241); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3243 = 5'ha == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_3242); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3244 = 5'hb == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_3243); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3245 = 5'hc == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_3244); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3246 = 5'hd == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_3245); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3247 = 5'he == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_3246); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3248 = 5'hf == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_3247); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3249 = 5'h10 == cnt[4:0] ? $signed(-32'sh10000) : $signed(_GEN_3248); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3250 = 5'h11 == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_3249); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3251 = 5'h12 == cnt[4:0] ? $signed(-32'shfb15) : $signed(_GEN_3250); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3252 = 5'h13 == cnt[4:0] ? $signed(-32'shf4fa) : $signed(_GEN_3251); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3253 = 5'h14 == cnt[4:0] ? $signed(-32'shec83) : $signed(_GEN_3252); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3254 = 5'h15 == cnt[4:0] ? $signed(-32'she1c6) : $signed(_GEN_3253); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3255 = 5'h16 == cnt[4:0] ? $signed(-32'shd4db) : $signed(_GEN_3254); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3256 = 5'h17 == cnt[4:0] ? $signed(-32'shc5e4) : $signed(_GEN_3255); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3257 = 5'h18 == cnt[4:0] ? $signed(-32'shb505) : $signed(_GEN_3256); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3258 = 5'h19 == cnt[4:0] ? $signed(-32'sha268) : $signed(_GEN_3257); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3259 = 5'h1a == cnt[4:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3258); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3260 = 5'h1b == cnt[4:0] ? $signed(-32'sh78ad) : $signed(_GEN_3259); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3261 = 5'h1c == cnt[4:0] ? $signed(-32'sh61f8) : $signed(_GEN_3260); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3262 = 5'h1d == cnt[4:0] ? $signed(-32'sh4a50) : $signed(_GEN_3261); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3263 = 5'h1e == cnt[4:0] ? $signed(-32'sh31f1) : $signed(_GEN_3262); // @[FFT.scala 52:18]
  reg [31:0] _T_849_re; // @[Reg.scala 15:16]
  reg [31:0] _T_849_im; // @[Reg.scala 15:16]
  reg [31:0] _T_850_re; // @[Reg.scala 15:16]
  reg [31:0] _T_850_im; // @[Reg.scala 15:16]
  reg [31:0] _T_851_re; // @[Reg.scala 15:16]
  reg [31:0] _T_851_im; // @[Reg.scala 15:16]
  reg [31:0] _T_852_re; // @[Reg.scala 15:16]
  reg [31:0] _T_852_im; // @[Reg.scala 15:16]
  reg [31:0] _T_853_re; // @[Reg.scala 15:16]
  reg [31:0] _T_853_im; // @[Reg.scala 15:16]
  reg [31:0] _T_854_re; // @[Reg.scala 15:16]
  reg [31:0] _T_854_im; // @[Reg.scala 15:16]
  reg [31:0] _T_855_re; // @[Reg.scala 15:16]
  reg [31:0] _T_855_im; // @[Reg.scala 15:16]
  reg [31:0] _T_856_re; // @[Reg.scala 15:16]
  reg [31:0] _T_856_im; // @[Reg.scala 15:16]
  reg [31:0] _T_857_re; // @[Reg.scala 15:16]
  reg [31:0] _T_857_im; // @[Reg.scala 15:16]
  reg [31:0] _T_858_re; // @[Reg.scala 15:16]
  reg [31:0] _T_858_im; // @[Reg.scala 15:16]
  reg [31:0] _T_859_re; // @[Reg.scala 15:16]
  reg [31:0] _T_859_im; // @[Reg.scala 15:16]
  reg [31:0] _T_860_re; // @[Reg.scala 15:16]
  reg [31:0] _T_860_im; // @[Reg.scala 15:16]
  reg [31:0] _T_861_re; // @[Reg.scala 15:16]
  reg [31:0] _T_861_im; // @[Reg.scala 15:16]
  reg [31:0] _T_862_re; // @[Reg.scala 15:16]
  reg [31:0] _T_862_im; // @[Reg.scala 15:16]
  reg [31:0] _T_863_re; // @[Reg.scala 15:16]
  reg [31:0] _T_863_im; // @[Reg.scala 15:16]
  reg [31:0] _T_864_re; // @[Reg.scala 15:16]
  reg [31:0] _T_864_im; // @[Reg.scala 15:16]
  reg [31:0] _T_865_re; // @[Reg.scala 15:16]
  reg [31:0] _T_865_im; // @[Reg.scala 15:16]
  reg [31:0] _T_866_re; // @[Reg.scala 15:16]
  reg [31:0] _T_866_im; // @[Reg.scala 15:16]
  reg [31:0] _T_867_re; // @[Reg.scala 15:16]
  reg [31:0] _T_867_im; // @[Reg.scala 15:16]
  reg [31:0] _T_868_re; // @[Reg.scala 15:16]
  reg [31:0] _T_868_im; // @[Reg.scala 15:16]
  reg [31:0] _T_869_re; // @[Reg.scala 15:16]
  reg [31:0] _T_869_im; // @[Reg.scala 15:16]
  reg [31:0] _T_870_re; // @[Reg.scala 15:16]
  reg [31:0] _T_870_im; // @[Reg.scala 15:16]
  reg [31:0] _T_871_re; // @[Reg.scala 15:16]
  reg [31:0] _T_871_im; // @[Reg.scala 15:16]
  reg [31:0] _T_872_re; // @[Reg.scala 15:16]
  reg [31:0] _T_872_im; // @[Reg.scala 15:16]
  reg [31:0] _T_873_re; // @[Reg.scala 15:16]
  reg [31:0] _T_873_im; // @[Reg.scala 15:16]
  reg [31:0] _T_874_re; // @[Reg.scala 15:16]
  reg [31:0] _T_874_im; // @[Reg.scala 15:16]
  reg [31:0] _T_875_re; // @[Reg.scala 15:16]
  reg [31:0] _T_875_im; // @[Reg.scala 15:16]
  reg [31:0] _T_876_re; // @[Reg.scala 15:16]
  reg [31:0] _T_876_im; // @[Reg.scala 15:16]
  reg [31:0] _T_877_re; // @[Reg.scala 15:16]
  reg [31:0] _T_877_im; // @[Reg.scala 15:16]
  reg [31:0] _T_878_re; // @[Reg.scala 15:16]
  reg [31:0] _T_878_im; // @[Reg.scala 15:16]
  reg [31:0] _T_879_re; // @[Reg.scala 15:16]
  reg [31:0] _T_879_im; // @[Reg.scala 15:16]
  reg [31:0] _T_880_re; // @[Reg.scala 15:16]
  reg [31:0] _T_880_im; // @[Reg.scala 15:16]
  reg [31:0] _T_882_re; // @[Reg.scala 15:16]
  reg [31:0] _T_882_im; // @[Reg.scala 15:16]
  reg [31:0] _T_883_re; // @[Reg.scala 15:16]
  reg [31:0] _T_883_im; // @[Reg.scala 15:16]
  reg [31:0] _T_884_re; // @[Reg.scala 15:16]
  reg [31:0] _T_884_im; // @[Reg.scala 15:16]
  reg [31:0] _T_885_re; // @[Reg.scala 15:16]
  reg [31:0] _T_885_im; // @[Reg.scala 15:16]
  reg [31:0] _T_886_re; // @[Reg.scala 15:16]
  reg [31:0] _T_886_im; // @[Reg.scala 15:16]
  reg [31:0] _T_887_re; // @[Reg.scala 15:16]
  reg [31:0] _T_887_im; // @[Reg.scala 15:16]
  reg [31:0] _T_888_re; // @[Reg.scala 15:16]
  reg [31:0] _T_888_im; // @[Reg.scala 15:16]
  reg [31:0] _T_889_re; // @[Reg.scala 15:16]
  reg [31:0] _T_889_im; // @[Reg.scala 15:16]
  reg [31:0] _T_890_re; // @[Reg.scala 15:16]
  reg [31:0] _T_890_im; // @[Reg.scala 15:16]
  reg [31:0] _T_891_re; // @[Reg.scala 15:16]
  reg [31:0] _T_891_im; // @[Reg.scala 15:16]
  reg [31:0] _T_892_re; // @[Reg.scala 15:16]
  reg [31:0] _T_892_im; // @[Reg.scala 15:16]
  reg [31:0] _T_893_re; // @[Reg.scala 15:16]
  reg [31:0] _T_893_im; // @[Reg.scala 15:16]
  reg [31:0] _T_894_re; // @[Reg.scala 15:16]
  reg [31:0] _T_894_im; // @[Reg.scala 15:16]
  reg [31:0] _T_895_re; // @[Reg.scala 15:16]
  reg [31:0] _T_895_im; // @[Reg.scala 15:16]
  reg [31:0] _T_896_re; // @[Reg.scala 15:16]
  reg [31:0] _T_896_im; // @[Reg.scala 15:16]
  reg [31:0] _T_897_re; // @[Reg.scala 15:16]
  reg [31:0] _T_897_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3362 = 4'h1 == cnt[3:0] ? $signed(32'shfb15) : $signed(32'sh10000); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3363 = 4'h2 == cnt[3:0] ? $signed(32'shec83) : $signed(_GEN_3362); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3364 = 4'h3 == cnt[3:0] ? $signed(32'shd4db) : $signed(_GEN_3363); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3365 = 4'h4 == cnt[3:0] ? $signed(32'shb505) : $signed(_GEN_3364); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3366 = 4'h5 == cnt[3:0] ? $signed(32'sh8e3a) : $signed(_GEN_3365); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3367 = 4'h6 == cnt[3:0] ? $signed(32'sh61f8) : $signed(_GEN_3366); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3368 = 4'h7 == cnt[3:0] ? $signed(32'sh31f1) : $signed(_GEN_3367); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3369 = 4'h8 == cnt[3:0] ? $signed(32'sh0) : $signed(_GEN_3368); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3370 = 4'h9 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_3369); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3371 = 4'ha == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_3370); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3372 = 4'hb == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3371); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3373 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_3372); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3374 = 4'hd == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_3373); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3375 = 4'he == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_3374); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3410 = 4'h1 == cnt[3:0] ? $signed(-32'sh31f1) : $signed(32'sh0); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3411 = 4'h2 == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_3410); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3412 = 4'h3 == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3411); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3413 = 4'h4 == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_3412); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3414 = 4'h5 == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_3413); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3415 = 4'h6 == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_3414); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3416 = 4'h7 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_3415); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3417 = 4'h8 == cnt[3:0] ? $signed(-32'sh10000) : $signed(_GEN_3416); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3418 = 4'h9 == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_3417); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3419 = 4'ha == cnt[3:0] ? $signed(-32'shec83) : $signed(_GEN_3418); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3420 = 4'hb == cnt[3:0] ? $signed(-32'shd4db) : $signed(_GEN_3419); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3421 = 4'hc == cnt[3:0] ? $signed(-32'shb505) : $signed(_GEN_3420); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3422 = 4'hd == cnt[3:0] ? $signed(-32'sh8e3a) : $signed(_GEN_3421); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3423 = 4'he == cnt[3:0] ? $signed(-32'sh61f8) : $signed(_GEN_3422); // @[FFT.scala 52:18]
  reg [31:0] _T_906_re; // @[Reg.scala 15:16]
  reg [31:0] _T_906_im; // @[Reg.scala 15:16]
  reg [31:0] _T_907_re; // @[Reg.scala 15:16]
  reg [31:0] _T_907_im; // @[Reg.scala 15:16]
  reg [31:0] _T_908_re; // @[Reg.scala 15:16]
  reg [31:0] _T_908_im; // @[Reg.scala 15:16]
  reg [31:0] _T_909_re; // @[Reg.scala 15:16]
  reg [31:0] _T_909_im; // @[Reg.scala 15:16]
  reg [31:0] _T_910_re; // @[Reg.scala 15:16]
  reg [31:0] _T_910_im; // @[Reg.scala 15:16]
  reg [31:0] _T_911_re; // @[Reg.scala 15:16]
  reg [31:0] _T_911_im; // @[Reg.scala 15:16]
  reg [31:0] _T_912_re; // @[Reg.scala 15:16]
  reg [31:0] _T_912_im; // @[Reg.scala 15:16]
  reg [31:0] _T_913_re; // @[Reg.scala 15:16]
  reg [31:0] _T_913_im; // @[Reg.scala 15:16]
  reg [31:0] _T_914_re; // @[Reg.scala 15:16]
  reg [31:0] _T_914_im; // @[Reg.scala 15:16]
  reg [31:0] _T_915_re; // @[Reg.scala 15:16]
  reg [31:0] _T_915_im; // @[Reg.scala 15:16]
  reg [31:0] _T_916_re; // @[Reg.scala 15:16]
  reg [31:0] _T_916_im; // @[Reg.scala 15:16]
  reg [31:0] _T_917_re; // @[Reg.scala 15:16]
  reg [31:0] _T_917_im; // @[Reg.scala 15:16]
  reg [31:0] _T_918_re; // @[Reg.scala 15:16]
  reg [31:0] _T_918_im; // @[Reg.scala 15:16]
  reg [31:0] _T_919_re; // @[Reg.scala 15:16]
  reg [31:0] _T_919_im; // @[Reg.scala 15:16]
  reg [31:0] _T_920_re; // @[Reg.scala 15:16]
  reg [31:0] _T_920_im; // @[Reg.scala 15:16]
  reg [31:0] _T_921_re; // @[Reg.scala 15:16]
  reg [31:0] _T_921_im; // @[Reg.scala 15:16]
  reg [31:0] _T_923_re; // @[Reg.scala 15:16]
  reg [31:0] _T_923_im; // @[Reg.scala 15:16]
  reg [31:0] _T_924_re; // @[Reg.scala 15:16]
  reg [31:0] _T_924_im; // @[Reg.scala 15:16]
  reg [31:0] _T_925_re; // @[Reg.scala 15:16]
  reg [31:0] _T_925_im; // @[Reg.scala 15:16]
  reg [31:0] _T_926_re; // @[Reg.scala 15:16]
  reg [31:0] _T_926_im; // @[Reg.scala 15:16]
  reg [31:0] _T_927_re; // @[Reg.scala 15:16]
  reg [31:0] _T_927_im; // @[Reg.scala 15:16]
  reg [31:0] _T_928_re; // @[Reg.scala 15:16]
  reg [31:0] _T_928_im; // @[Reg.scala 15:16]
  reg [31:0] _T_929_re; // @[Reg.scala 15:16]
  reg [31:0] _T_929_im; // @[Reg.scala 15:16]
  reg [31:0] _T_930_re; // @[Reg.scala 15:16]
  reg [31:0] _T_930_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3474 = 3'h1 == cnt[2:0] ? $signed(32'shec83) : $signed(32'sh10000); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3475 = 3'h2 == cnt[2:0] ? $signed(32'shb505) : $signed(_GEN_3474); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3476 = 3'h3 == cnt[2:0] ? $signed(32'sh61f8) : $signed(_GEN_3475); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3477 = 3'h4 == cnt[2:0] ? $signed(32'sh0) : $signed(_GEN_3476); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3478 = 3'h5 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_3477); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3479 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_3478); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3498 = 3'h1 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(32'sh0); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3499 = 3'h2 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_3498); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3500 = 3'h3 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_3499); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3501 = 3'h4 == cnt[2:0] ? $signed(-32'sh10000) : $signed(_GEN_3500); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3502 = 3'h5 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_3501); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3503 = 3'h6 == cnt[2:0] ? $signed(-32'shb505) : $signed(_GEN_3502); // @[FFT.scala 52:18]
  reg [31:0] _T_939_re; // @[Reg.scala 15:16]
  reg [31:0] _T_939_im; // @[Reg.scala 15:16]
  reg [31:0] _T_940_re; // @[Reg.scala 15:16]
  reg [31:0] _T_940_im; // @[Reg.scala 15:16]
  reg [31:0] _T_941_re; // @[Reg.scala 15:16]
  reg [31:0] _T_941_im; // @[Reg.scala 15:16]
  reg [31:0] _T_942_re; // @[Reg.scala 15:16]
  reg [31:0] _T_942_im; // @[Reg.scala 15:16]
  reg [31:0] _T_943_re; // @[Reg.scala 15:16]
  reg [31:0] _T_943_im; // @[Reg.scala 15:16]
  reg [31:0] _T_944_re; // @[Reg.scala 15:16]
  reg [31:0] _T_944_im; // @[Reg.scala 15:16]
  reg [31:0] _T_945_re; // @[Reg.scala 15:16]
  reg [31:0] _T_945_im; // @[Reg.scala 15:16]
  reg [31:0] _T_946_re; // @[Reg.scala 15:16]
  reg [31:0] _T_946_im; // @[Reg.scala 15:16]
  reg [31:0] _T_948_re; // @[Reg.scala 15:16]
  reg [31:0] _T_948_im; // @[Reg.scala 15:16]
  reg [31:0] _T_949_re; // @[Reg.scala 15:16]
  reg [31:0] _T_949_im; // @[Reg.scala 15:16]
  reg [31:0] _T_950_re; // @[Reg.scala 15:16]
  reg [31:0] _T_950_im; // @[Reg.scala 15:16]
  reg [31:0] _T_951_re; // @[Reg.scala 15:16]
  reg [31:0] _T_951_im; // @[Reg.scala 15:16]
  wire [31:0] _GEN_3530 = 2'h1 == cnt[1:0] ? $signed(32'shb505) : $signed(32'sh10000); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3531 = 2'h2 == cnt[1:0] ? $signed(32'sh0) : $signed(_GEN_3530); // @[FFT.scala 51:18]
  wire [31:0] _GEN_3542 = 2'h1 == cnt[1:0] ? $signed(-32'shb505) : $signed(32'sh0); // @[FFT.scala 52:18]
  wire [31:0] _GEN_3543 = 2'h2 == cnt[1:0] ? $signed(-32'sh10000) : $signed(_GEN_3542); // @[FFT.scala 52:18]
  reg [31:0] _T_960_re; // @[Reg.scala 15:16]
  reg [31:0] _T_960_im; // @[Reg.scala 15:16]
  reg [31:0] _T_961_re; // @[Reg.scala 15:16]
  reg [31:0] _T_961_im; // @[Reg.scala 15:16]
  reg [31:0] _T_962_re; // @[Reg.scala 15:16]
  reg [31:0] _T_962_im; // @[Reg.scala 15:16]
  reg [31:0] _T_963_re; // @[Reg.scala 15:16]
  reg [31:0] _T_963_im; // @[Reg.scala 15:16]
  reg [31:0] _T_965_re; // @[Reg.scala 15:16]
  reg [31:0] _T_965_im; // @[Reg.scala 15:16]
  reg [31:0] _T_966_re; // @[Reg.scala 15:16]
  reg [31:0] _T_966_im; // @[Reg.scala 15:16]
  reg [31:0] _T_975_re; // @[Reg.scala 15:16]
  reg [31:0] _T_975_im; // @[Reg.scala 15:16]
  reg [31:0] _T_976_re; // @[Reg.scala 15:16]
  reg [31:0] _T_976_im; // @[Reg.scala 15:16]
  reg [31:0] _T_978_re; // @[Reg.scala 15:16]
  reg [31:0] _T_978_im; // @[Reg.scala 15:16]
  reg [31:0] out1D1_re; // @[FFT.scala 82:23]
  reg [31:0] out1D1_im; // @[FFT.scala 82:23]
  reg [31:0] _T_985_re; // @[FFT.scala 88:22]
  reg [31:0] _T_985_im; // @[FFT.scala 88:22]
  reg [31:0] _T_986_re; // @[FFT.scala 89:22]
  reg [31:0] _T_986_im; // @[FFT.scala 89:22]
  reg  _T_987; // @[Reg.scala 15:16]
  reg  _T_988; // @[Reg.scala 15:16]
  reg  _T_989; // @[Reg.scala 15:16]
  reg  _T_990; // @[Reg.scala 15:16]
  reg  _T_991; // @[Reg.scala 15:16]
  reg  _T_992; // @[Reg.scala 15:16]
  reg  _T_993; // @[Reg.scala 15:16]
  reg  _T_994; // @[Reg.scala 15:16]
  reg  _T_995; // @[Reg.scala 15:16]
  reg  _T_996; // @[Reg.scala 15:16]
  reg  _T_997; // @[Reg.scala 15:16]
  reg  _T_998; // @[Reg.scala 15:16]
  reg  _T_999; // @[Reg.scala 15:16]
  reg  _T_1000; // @[Reg.scala 15:16]
  reg  _T_1001; // @[Reg.scala 15:16]
  reg  _T_1002; // @[Reg.scala 15:16]
  reg  _T_1003; // @[Reg.scala 15:16]
  reg  _T_1004; // @[Reg.scala 15:16]
  reg  _T_1005; // @[Reg.scala 15:16]
  reg  _T_1006; // @[Reg.scala 15:16]
  reg  _T_1007; // @[Reg.scala 15:16]
  reg  _T_1008; // @[Reg.scala 15:16]
  reg  _T_1009; // @[Reg.scala 15:16]
  reg  _T_1010; // @[Reg.scala 15:16]
  reg  _T_1011; // @[Reg.scala 15:16]
  reg  _T_1012; // @[Reg.scala 15:16]
  reg  _T_1013; // @[Reg.scala 15:16]
  reg  _T_1014; // @[Reg.scala 15:16]
  reg  _T_1015; // @[Reg.scala 15:16]
  reg  _T_1016; // @[Reg.scala 15:16]
  reg  _T_1017; // @[Reg.scala 15:16]
  reg  _T_1018; // @[Reg.scala 15:16]
  reg  _T_1019; // @[Reg.scala 15:16]
  reg  _T_1020; // @[Reg.scala 15:16]
  reg  _T_1021; // @[Reg.scala 15:16]
  reg  _T_1022; // @[Reg.scala 15:16]
  reg  _T_1023; // @[Reg.scala 15:16]
  reg  _T_1024; // @[Reg.scala 15:16]
  reg  _T_1025; // @[Reg.scala 15:16]
  reg  _T_1026; // @[Reg.scala 15:16]
  reg  _T_1027; // @[Reg.scala 15:16]
  reg  _T_1028; // @[Reg.scala 15:16]
  reg  _T_1029; // @[Reg.scala 15:16]
  reg  _T_1030; // @[Reg.scala 15:16]
  reg  _T_1031; // @[Reg.scala 15:16]
  reg  _T_1032; // @[Reg.scala 15:16]
  reg  _T_1033; // @[Reg.scala 15:16]
  reg  _T_1034; // @[Reg.scala 15:16]
  reg  _T_1035; // @[Reg.scala 15:16]
  reg  _T_1036; // @[Reg.scala 15:16]
  reg  _T_1037; // @[Reg.scala 15:16]
  reg  _T_1038; // @[Reg.scala 15:16]
  reg  _T_1039; // @[Reg.scala 15:16]
  reg  _T_1040; // @[Reg.scala 15:16]
  reg  _T_1041; // @[Reg.scala 15:16]
  reg  _T_1042; // @[Reg.scala 15:16]
  reg  _T_1043; // @[Reg.scala 15:16]
  reg  _T_1044; // @[Reg.scala 15:16]
  reg  _T_1045; // @[Reg.scala 15:16]
  reg  _T_1046; // @[Reg.scala 15:16]
  reg  _T_1047; // @[Reg.scala 15:16]
  reg  _T_1048; // @[Reg.scala 15:16]
  reg  _T_1049; // @[Reg.scala 15:16]
  reg  _T_1050; // @[Reg.scala 15:16]
  reg  _T_1051; // @[Reg.scala 15:16]
  reg  _T_1052; // @[Reg.scala 15:16]
  reg  _T_1053; // @[Reg.scala 15:16]
  reg  _T_1054; // @[Reg.scala 15:16]
  reg  _T_1055; // @[Reg.scala 15:16]
  reg  _T_1056; // @[Reg.scala 15:16]
  reg  _T_1057; // @[Reg.scala 15:16]
  reg  _T_1058; // @[Reg.scala 15:16]
  reg  _T_1059; // @[Reg.scala 15:16]
  reg  _T_1060; // @[Reg.scala 15:16]
  reg  _T_1061; // @[Reg.scala 15:16]
  reg  _T_1062; // @[Reg.scala 15:16]
  reg  _T_1063; // @[Reg.scala 15:16]
  reg  _T_1064; // @[Reg.scala 15:16]
  reg  _T_1065; // @[Reg.scala 15:16]
  reg  _T_1066; // @[Reg.scala 15:16]
  reg  _T_1067; // @[Reg.scala 15:16]
  reg  _T_1068; // @[Reg.scala 15:16]
  reg  _T_1069; // @[Reg.scala 15:16]
  reg  _T_1070; // @[Reg.scala 15:16]
  reg  _T_1071; // @[Reg.scala 15:16]
  reg  _T_1072; // @[Reg.scala 15:16]
  reg  _T_1073; // @[Reg.scala 15:16]
  reg  _T_1074; // @[Reg.scala 15:16]
  reg  _T_1075; // @[Reg.scala 15:16]
  reg  _T_1076; // @[Reg.scala 15:16]
  reg  _T_1077; // @[Reg.scala 15:16]
  reg  _T_1078; // @[Reg.scala 15:16]
  reg  _T_1079; // @[Reg.scala 15:16]
  reg  _T_1080; // @[Reg.scala 15:16]
  reg  _T_1081; // @[Reg.scala 15:16]
  reg  _T_1082; // @[Reg.scala 15:16]
  reg  _T_1083; // @[Reg.scala 15:16]
  reg  _T_1084; // @[Reg.scala 15:16]
  reg  _T_1085; // @[Reg.scala 15:16]
  reg  _T_1086; // @[Reg.scala 15:16]
  reg  _T_1087; // @[Reg.scala 15:16]
  reg  _T_1088; // @[Reg.scala 15:16]
  reg  _T_1089; // @[Reg.scala 15:16]
  reg  _T_1090; // @[Reg.scala 15:16]
  reg  _T_1091; // @[Reg.scala 15:16]
  reg  _T_1092; // @[Reg.scala 15:16]
  reg  _T_1093; // @[Reg.scala 15:16]
  reg  _T_1094; // @[Reg.scala 15:16]
  reg  _T_1095; // @[Reg.scala 15:16]
  reg  _T_1096; // @[Reg.scala 15:16]
  reg  _T_1097; // @[Reg.scala 15:16]
  reg  _T_1098; // @[Reg.scala 15:16]
  reg  _T_1099; // @[Reg.scala 15:16]
  reg  _T_1100; // @[Reg.scala 15:16]
  reg  _T_1101; // @[Reg.scala 15:16]
  reg  _T_1102; // @[Reg.scala 15:16]
  reg  _T_1103; // @[Reg.scala 15:16]
  reg  _T_1104; // @[Reg.scala 15:16]
  reg  _T_1105; // @[Reg.scala 15:16]
  reg  _T_1106; // @[Reg.scala 15:16]
  reg  _T_1107; // @[Reg.scala 15:16]
  reg  _T_1108; // @[Reg.scala 15:16]
  reg  _T_1109; // @[Reg.scala 15:16]
  reg  _T_1110; // @[Reg.scala 15:16]
  reg  _T_1111; // @[Reg.scala 15:16]
  reg  _T_1112; // @[Reg.scala 15:16]
  reg  _T_1113; // @[Reg.scala 15:16]
  reg  _T_1114; // @[Reg.scala 15:16]
  reg  _T_1115; // @[Reg.scala 15:16]
  reg  _T_1116; // @[Reg.scala 15:16]
  reg  _T_1117; // @[Reg.scala 15:16]
  reg  _T_1118; // @[Reg.scala 15:16]
  reg  _T_1119; // @[Reg.scala 15:16]
  reg  _T_1120; // @[Reg.scala 15:16]
  reg  _T_1121; // @[Reg.scala 15:16]
  reg  _T_1122; // @[Reg.scala 15:16]
  reg  _T_1123; // @[Reg.scala 15:16]
  reg  _T_1124; // @[Reg.scala 15:16]
  reg  _T_1125; // @[Reg.scala 15:16]
  reg  _T_1126; // @[Reg.scala 15:16]
  reg  _T_1127; // @[Reg.scala 15:16]
  reg  _T_1128; // @[Reg.scala 15:16]
  reg  _T_1129; // @[Reg.scala 15:16]
  reg  _T_1130; // @[Reg.scala 15:16]
  reg  _T_1131; // @[Reg.scala 15:16]
  reg  _T_1132; // @[Reg.scala 15:16]
  reg  _T_1133; // @[Reg.scala 15:16]
  reg  _T_1134; // @[Reg.scala 15:16]
  reg  _T_1135; // @[Reg.scala 15:16]
  reg  _T_1136; // @[Reg.scala 15:16]
  reg  _T_1137; // @[Reg.scala 15:16]
  reg  _T_1138; // @[Reg.scala 15:16]
  reg  _T_1139; // @[Reg.scala 15:16]
  reg  _T_1140; // @[Reg.scala 15:16]
  reg  _T_1141; // @[Reg.scala 15:16]
  reg  _T_1142; // @[Reg.scala 15:16]
  reg  _T_1143; // @[Reg.scala 15:16]
  reg  _T_1144; // @[Reg.scala 15:16]
  reg  _T_1145; // @[Reg.scala 15:16]
  reg  _T_1146; // @[Reg.scala 15:16]
  reg  _T_1147; // @[Reg.scala 15:16]
  reg  _T_1148; // @[Reg.scala 15:16]
  reg  _T_1149; // @[Reg.scala 15:16]
  reg  _T_1150; // @[Reg.scala 15:16]
  reg  _T_1151; // @[Reg.scala 15:16]
  reg  _T_1152; // @[Reg.scala 15:16]
  reg  _T_1153; // @[Reg.scala 15:16]
  reg  _T_1154; // @[Reg.scala 15:16]
  reg  _T_1155; // @[Reg.scala 15:16]
  reg  _T_1156; // @[Reg.scala 15:16]
  reg  _T_1157; // @[Reg.scala 15:16]
  reg  _T_1158; // @[Reg.scala 15:16]
  reg  _T_1159; // @[Reg.scala 15:16]
  reg  _T_1160; // @[Reg.scala 15:16]
  reg  _T_1161; // @[Reg.scala 15:16]
  reg  _T_1162; // @[Reg.scala 15:16]
  reg  _T_1163; // @[Reg.scala 15:16]
  reg  _T_1164; // @[Reg.scala 15:16]
  reg  _T_1165; // @[Reg.scala 15:16]
  reg  _T_1166; // @[Reg.scala 15:16]
  reg  _T_1167; // @[Reg.scala 15:16]
  reg  _T_1168; // @[Reg.scala 15:16]
  reg  _T_1169; // @[Reg.scala 15:16]
  reg  _T_1170; // @[Reg.scala 15:16]
  reg  _T_1171; // @[Reg.scala 15:16]
  reg  _T_1172; // @[Reg.scala 15:16]
  reg  _T_1173; // @[Reg.scala 15:16]
  reg  _T_1174; // @[Reg.scala 15:16]
  reg  _T_1175; // @[Reg.scala 15:16]
  reg  _T_1176; // @[Reg.scala 15:16]
  reg  _T_1177; // @[Reg.scala 15:16]
  reg  _T_1178; // @[Reg.scala 15:16]
  reg  _T_1179; // @[Reg.scala 15:16]
  reg  _T_1180; // @[Reg.scala 15:16]
  reg  _T_1181; // @[Reg.scala 15:16]
  reg  _T_1182; // @[Reg.scala 15:16]
  reg  _T_1183; // @[Reg.scala 15:16]
  reg  _T_1184; // @[Reg.scala 15:16]
  reg  _T_1185; // @[Reg.scala 15:16]
  reg  _T_1186; // @[Reg.scala 15:16]
  reg  _T_1187; // @[Reg.scala 15:16]
  reg  _T_1188; // @[Reg.scala 15:16]
  reg  _T_1189; // @[Reg.scala 15:16]
  reg  _T_1190; // @[Reg.scala 15:16]
  reg  _T_1191; // @[Reg.scala 15:16]
  reg  _T_1192; // @[Reg.scala 15:16]
  reg  _T_1193; // @[Reg.scala 15:16]
  reg  _T_1194; // @[Reg.scala 15:16]
  reg  _T_1195; // @[Reg.scala 15:16]
  reg  _T_1196; // @[Reg.scala 15:16]
  reg  _T_1197; // @[Reg.scala 15:16]
  reg  _T_1198; // @[Reg.scala 15:16]
  reg  _T_1199; // @[Reg.scala 15:16]
  reg  _T_1200; // @[Reg.scala 15:16]
  reg  _T_1201; // @[Reg.scala 15:16]
  reg  _T_1202; // @[Reg.scala 15:16]
  reg  _T_1203; // @[Reg.scala 15:16]
  reg  _T_1204; // @[Reg.scala 15:16]
  reg  _T_1205; // @[Reg.scala 15:16]
  reg  _T_1206; // @[Reg.scala 15:16]
  reg  _T_1207; // @[Reg.scala 15:16]
  reg  _T_1208; // @[Reg.scala 15:16]
  reg  _T_1209; // @[Reg.scala 15:16]
  reg  _T_1210; // @[Reg.scala 15:16]
  reg  _T_1211; // @[Reg.scala 15:16]
  reg  _T_1212; // @[Reg.scala 15:16]
  reg  _T_1213; // @[Reg.scala 15:16]
  reg  _T_1214; // @[Reg.scala 15:16]
  reg  _T_1215; // @[Reg.scala 15:16]
  reg  _T_1216; // @[Reg.scala 15:16]
  reg  _T_1217; // @[Reg.scala 15:16]
  reg  _T_1218; // @[Reg.scala 15:16]
  reg  _T_1219; // @[Reg.scala 15:16]
  reg  _T_1220; // @[Reg.scala 15:16]
  reg  _T_1221; // @[Reg.scala 15:16]
  reg  _T_1222; // @[Reg.scala 15:16]
  reg  _T_1223; // @[Reg.scala 15:16]
  reg  _T_1224; // @[Reg.scala 15:16]
  reg  _T_1225; // @[Reg.scala 15:16]
  reg  _T_1226; // @[Reg.scala 15:16]
  reg  _T_1227; // @[Reg.scala 15:16]
  reg  _T_1228; // @[Reg.scala 15:16]
  reg  _T_1229; // @[Reg.scala 15:16]
  reg  _T_1230; // @[Reg.scala 15:16]
  reg  _T_1231; // @[Reg.scala 15:16]
  reg  _T_1232; // @[Reg.scala 15:16]
  reg  _T_1233; // @[Reg.scala 15:16]
  reg  _T_1234; // @[Reg.scala 15:16]
  reg  _T_1235; // @[Reg.scala 15:16]
  reg  _T_1236; // @[Reg.scala 15:16]
  reg  _T_1237; // @[Reg.scala 15:16]
  reg  _T_1238; // @[Reg.scala 15:16]
  reg  _T_1239; // @[Reg.scala 15:16]
  reg  _T_1240; // @[Reg.scala 15:16]
  reg  _T_1241; // @[Reg.scala 15:16]
  reg  _T_1242; // @[Reg.scala 15:16]
  reg  _T_1243; // @[Reg.scala 15:16]
  reg  _T_1244; // @[Reg.scala 15:16]
  reg  _T_1245; // @[Reg.scala 15:16]
  reg  _T_1246; // @[Reg.scala 15:16]
  reg  _T_1247; // @[Reg.scala 15:16]
  reg  _T_1248; // @[Reg.scala 15:16]
  reg  _T_1249; // @[Reg.scala 15:16]
  reg  _T_1250; // @[Reg.scala 15:16]
  reg  _T_1251; // @[Reg.scala 15:16]
  reg  _T_1252; // @[Reg.scala 15:16]
  reg  _T_1253; // @[Reg.scala 15:16]
  reg  _T_1254; // @[Reg.scala 15:16]
  reg  _T_1255; // @[Reg.scala 15:16]
  reg  _T_1256; // @[Reg.scala 15:16]
  reg  _T_1257; // @[Reg.scala 15:16]
  reg  _T_1258; // @[Reg.scala 15:16]
  reg  _T_1259; // @[Reg.scala 15:16]
  reg  _T_1260; // @[Reg.scala 15:16]
  reg  _T_1261; // @[Reg.scala 15:16]
  reg  _T_1262; // @[Reg.scala 15:16]
  reg  _T_1263; // @[Reg.scala 15:16]
  reg  _T_1264; // @[Reg.scala 15:16]
  reg  _T_1265; // @[Reg.scala 15:16]
  reg  _T_1266; // @[Reg.scala 15:16]
  reg  _T_1267; // @[Reg.scala 15:16]
  reg  _T_1268; // @[Reg.scala 15:16]
  reg  _T_1269; // @[Reg.scala 15:16]
  reg  _T_1270; // @[Reg.scala 15:16]
  reg  _T_1271; // @[Reg.scala 15:16]
  reg  _T_1272; // @[Reg.scala 15:16]
  reg  _T_1273; // @[Reg.scala 15:16]
  reg  _T_1274; // @[Reg.scala 15:16]
  reg  _T_1275; // @[Reg.scala 15:16]
  reg  _T_1276; // @[Reg.scala 15:16]
  reg  _T_1277; // @[Reg.scala 15:16]
  reg  _T_1278; // @[Reg.scala 15:16]
  reg  _T_1279; // @[Reg.scala 15:16]
  reg  _T_1280; // @[Reg.scala 15:16]
  reg  _T_1281; // @[Reg.scala 15:16]
  reg  _T_1282; // @[Reg.scala 15:16]
  reg  _T_1283; // @[Reg.scala 15:16]
  reg  _T_1284; // @[Reg.scala 15:16]
  reg  _T_1285; // @[Reg.scala 15:16]
  reg  _T_1286; // @[Reg.scala 15:16]
  reg  _T_1287; // @[Reg.scala 15:16]
  reg  _T_1288; // @[Reg.scala 15:16]
  reg  _T_1289; // @[Reg.scala 15:16]
  reg  _T_1290; // @[Reg.scala 15:16]
  reg  _T_1291; // @[Reg.scala 15:16]
  reg  _T_1292; // @[Reg.scala 15:16]
  reg  _T_1293; // @[Reg.scala 15:16]
  reg  _T_1294; // @[Reg.scala 15:16]
  reg  _T_1295; // @[Reg.scala 15:16]
  reg  _T_1296; // @[Reg.scala 15:16]
  reg  _T_1297; // @[Reg.scala 15:16]
  reg  _T_1298; // @[Reg.scala 15:16]
  reg  _T_1299; // @[Reg.scala 15:16]
  reg  _T_1300; // @[Reg.scala 15:16]
  reg  _T_1301; // @[Reg.scala 15:16]
  reg  _T_1302; // @[Reg.scala 15:16]
  reg  _T_1303; // @[Reg.scala 15:16]
  reg  _T_1304; // @[Reg.scala 15:16]
  reg  _T_1305; // @[Reg.scala 15:16]
  reg  _T_1306; // @[Reg.scala 15:16]
  reg  _T_1307; // @[Reg.scala 15:16]
  reg  _T_1308; // @[Reg.scala 15:16]
  reg  _T_1309; // @[Reg.scala 15:16]
  reg  _T_1310; // @[Reg.scala 15:16]
  reg  _T_1311; // @[Reg.scala 15:16]
  reg  _T_1312; // @[Reg.scala 15:16]
  reg  _T_1313; // @[Reg.scala 15:16]
  reg  _T_1314; // @[Reg.scala 15:16]
  reg  _T_1315; // @[Reg.scala 15:16]
  reg  _T_1316; // @[Reg.scala 15:16]
  reg  _T_1317; // @[Reg.scala 15:16]
  reg  _T_1318; // @[Reg.scala 15:16]
  reg  _T_1319; // @[Reg.scala 15:16]
  reg  _T_1320; // @[Reg.scala 15:16]
  reg  _T_1321; // @[Reg.scala 15:16]
  reg  _T_1322; // @[Reg.scala 15:16]
  reg  _T_1323; // @[Reg.scala 15:16]
  reg  _T_1324; // @[Reg.scala 15:16]
  reg  _T_1325; // @[Reg.scala 15:16]
  reg  _T_1326; // @[Reg.scala 15:16]
  reg  _T_1327; // @[Reg.scala 15:16]
  reg  _T_1328; // @[Reg.scala 15:16]
  reg  _T_1329; // @[Reg.scala 15:16]
  reg  _T_1330; // @[Reg.scala 15:16]
  reg  _T_1331; // @[Reg.scala 15:16]
  reg  _T_1332; // @[Reg.scala 15:16]
  reg  _T_1333; // @[Reg.scala 15:16]
  reg  _T_1334; // @[Reg.scala 15:16]
  reg  _T_1335; // @[Reg.scala 15:16]
  reg  _T_1336; // @[Reg.scala 15:16]
  reg  _T_1337; // @[Reg.scala 15:16]
  reg  _T_1338; // @[Reg.scala 15:16]
  reg  _T_1339; // @[Reg.scala 15:16]
  reg  _T_1340; // @[Reg.scala 15:16]
  reg  _T_1341; // @[Reg.scala 15:16]
  reg  _T_1342; // @[Reg.scala 15:16]
  reg  _T_1343; // @[Reg.scala 15:16]
  reg  _T_1344; // @[Reg.scala 15:16]
  reg  _T_1345; // @[Reg.scala 15:16]
  reg  _T_1346; // @[Reg.scala 15:16]
  reg  _T_1347; // @[Reg.scala 15:16]
  reg  _T_1348; // @[Reg.scala 15:16]
  reg  _T_1349; // @[Reg.scala 15:16]
  reg  _T_1350; // @[Reg.scala 15:16]
  reg  _T_1351; // @[Reg.scala 15:16]
  reg  _T_1352; // @[Reg.scala 15:16]
  reg  _T_1353; // @[Reg.scala 15:16]
  reg  _T_1354; // @[Reg.scala 15:16]
  reg  _T_1355; // @[Reg.scala 15:16]
  reg  _T_1356; // @[Reg.scala 15:16]
  reg  _T_1357; // @[Reg.scala 15:16]
  reg  _T_1358; // @[Reg.scala 15:16]
  reg  _T_1359; // @[Reg.scala 15:16]
  reg  _T_1360; // @[Reg.scala 15:16]
  reg  _T_1361; // @[Reg.scala 15:16]
  reg  _T_1362; // @[Reg.scala 15:16]
  reg  _T_1363; // @[Reg.scala 15:16]
  reg  _T_1364; // @[Reg.scala 15:16]
  reg  _T_1365; // @[Reg.scala 15:16]
  reg  _T_1366; // @[Reg.scala 15:16]
  reg  _T_1367; // @[Reg.scala 15:16]
  reg  _T_1368; // @[Reg.scala 15:16]
  reg  _T_1369; // @[Reg.scala 15:16]
  reg  _T_1370; // @[Reg.scala 15:16]
  reg  _T_1371; // @[Reg.scala 15:16]
  reg  _T_1372; // @[Reg.scala 15:16]
  reg  _T_1373; // @[Reg.scala 15:16]
  reg  _T_1374; // @[Reg.scala 15:16]
  reg  _T_1375; // @[Reg.scala 15:16]
  reg  _T_1376; // @[Reg.scala 15:16]
  reg  _T_1377; // @[Reg.scala 15:16]
  reg  _T_1378; // @[Reg.scala 15:16]
  reg  _T_1379; // @[Reg.scala 15:16]
  reg  _T_1380; // @[Reg.scala 15:16]
  reg  _T_1381; // @[Reg.scala 15:16]
  reg  _T_1382; // @[Reg.scala 15:16]
  reg  _T_1383; // @[Reg.scala 15:16]
  reg  _T_1384; // @[Reg.scala 15:16]
  reg  _T_1385; // @[Reg.scala 15:16]
  reg  _T_1386; // @[Reg.scala 15:16]
  reg  _T_1387; // @[Reg.scala 15:16]
  reg  _T_1388; // @[Reg.scala 15:16]
  reg  _T_1389; // @[Reg.scala 15:16]
  reg  _T_1390; // @[Reg.scala 15:16]
  reg  _T_1391; // @[Reg.scala 15:16]
  reg  _T_1392; // @[Reg.scala 15:16]
  reg  _T_1393; // @[Reg.scala 15:16]
  reg  _T_1394; // @[Reg.scala 15:16]
  reg  _T_1395; // @[Reg.scala 15:16]
  reg  _T_1396; // @[Reg.scala 15:16]
  reg  _T_1397; // @[Reg.scala 15:16]
  reg  _T_1398; // @[Reg.scala 15:16]
  reg  _T_1399; // @[Reg.scala 15:16]
  reg  _T_1400; // @[Reg.scala 15:16]
  reg  _T_1401; // @[Reg.scala 15:16]
  reg  _T_1402; // @[Reg.scala 15:16]
  reg  _T_1403; // @[Reg.scala 15:16]
  reg  _T_1404; // @[Reg.scala 15:16]
  reg  _T_1405; // @[Reg.scala 15:16]
  reg  _T_1406; // @[Reg.scala 15:16]
  reg  _T_1407; // @[Reg.scala 15:16]
  reg  _T_1408; // @[Reg.scala 15:16]
  reg  _T_1409; // @[Reg.scala 15:16]
  reg  _T_1410; // @[Reg.scala 15:16]
  reg  _T_1411; // @[Reg.scala 15:16]
  reg  _T_1412; // @[Reg.scala 15:16]
  reg  _T_1413; // @[Reg.scala 15:16]
  reg  _T_1414; // @[Reg.scala 15:16]
  reg  _T_1415; // @[Reg.scala 15:16]
  reg  _T_1416; // @[Reg.scala 15:16]
  reg  _T_1417; // @[Reg.scala 15:16]
  reg  _T_1418; // @[Reg.scala 15:16]
  reg  _T_1419; // @[Reg.scala 15:16]
  reg  _T_1420; // @[Reg.scala 15:16]
  reg  _T_1421; // @[Reg.scala 15:16]
  reg  _T_1422; // @[Reg.scala 15:16]
  reg  _T_1423; // @[Reg.scala 15:16]
  reg  _T_1424; // @[Reg.scala 15:16]
  reg  _T_1425; // @[Reg.scala 15:16]
  reg  _T_1426; // @[Reg.scala 15:16]
  reg  _T_1427; // @[Reg.scala 15:16]
  reg  _T_1428; // @[Reg.scala 15:16]
  reg  _T_1429; // @[Reg.scala 15:16]
  reg  _T_1430; // @[Reg.scala 15:16]
  reg  _T_1431; // @[Reg.scala 15:16]
  reg  _T_1432; // @[Reg.scala 15:16]
  reg  _T_1433; // @[Reg.scala 15:16]
  reg  _T_1434; // @[Reg.scala 15:16]
  reg  _T_1435; // @[Reg.scala 15:16]
  reg  _T_1436; // @[Reg.scala 15:16]
  reg  _T_1437; // @[Reg.scala 15:16]
  reg  _T_1438; // @[Reg.scala 15:16]
  reg  _T_1439; // @[Reg.scala 15:16]
  reg  _T_1440; // @[Reg.scala 15:16]
  reg  _T_1441; // @[Reg.scala 15:16]
  reg  _T_1442; // @[Reg.scala 15:16]
  reg  _T_1443; // @[Reg.scala 15:16]
  reg  _T_1444; // @[Reg.scala 15:16]
  reg  _T_1445; // @[Reg.scala 15:16]
  reg  _T_1446; // @[Reg.scala 15:16]
  reg  _T_1447; // @[Reg.scala 15:16]
  reg  _T_1448; // @[Reg.scala 15:16]
  reg  _T_1449; // @[Reg.scala 15:16]
  reg  _T_1450; // @[Reg.scala 15:16]
  reg  _T_1451; // @[Reg.scala 15:16]
  reg  _T_1452; // @[Reg.scala 15:16]
  reg  _T_1453; // @[Reg.scala 15:16]
  reg  _T_1454; // @[Reg.scala 15:16]
  reg  _T_1455; // @[Reg.scala 15:16]
  reg  _T_1456; // @[Reg.scala 15:16]
  reg  _T_1457; // @[Reg.scala 15:16]
  reg  _T_1458; // @[Reg.scala 15:16]
  reg  _T_1459; // @[Reg.scala 15:16]
  reg  _T_1460; // @[Reg.scala 15:16]
  reg  _T_1461; // @[Reg.scala 15:16]
  reg  _T_1462; // @[Reg.scala 15:16]
  reg  _T_1463; // @[Reg.scala 15:16]
  reg  _T_1464; // @[Reg.scala 15:16]
  reg  _T_1465; // @[Reg.scala 15:16]
  reg  _T_1466; // @[Reg.scala 15:16]
  reg  _T_1467; // @[Reg.scala 15:16]
  reg  _T_1468; // @[Reg.scala 15:16]
  reg  _T_1469; // @[Reg.scala 15:16]
  reg  _T_1470; // @[Reg.scala 15:16]
  reg  _T_1471; // @[Reg.scala 15:16]
  reg  _T_1472; // @[Reg.scala 15:16]
  reg  _T_1473; // @[Reg.scala 15:16]
  reg  _T_1474; // @[Reg.scala 15:16]
  reg  _T_1475; // @[Reg.scala 15:16]
  reg  _T_1476; // @[Reg.scala 15:16]
  reg  _T_1477; // @[Reg.scala 15:16]
  reg  _T_1478; // @[Reg.scala 15:16]
  reg  _T_1479; // @[Reg.scala 15:16]
  reg  _T_1480; // @[Reg.scala 15:16]
  reg  _T_1481; // @[Reg.scala 15:16]
  reg  _T_1482; // @[Reg.scala 15:16]
  reg  _T_1483; // @[Reg.scala 15:16]
  reg  _T_1484; // @[Reg.scala 15:16]
  reg  _T_1485; // @[Reg.scala 15:16]
  reg  _T_1486; // @[Reg.scala 15:16]
  reg  _T_1487; // @[Reg.scala 15:16]
  reg  _T_1488; // @[Reg.scala 15:16]
  reg  _T_1489; // @[Reg.scala 15:16]
  reg  _T_1490; // @[Reg.scala 15:16]
  reg  _T_1491; // @[Reg.scala 15:16]
  reg  _T_1492; // @[Reg.scala 15:16]
  reg  _T_1493; // @[Reg.scala 15:16]
  reg  _T_1494; // @[Reg.scala 15:16]
  reg  _T_1495; // @[Reg.scala 15:16]
  reg  _T_1496; // @[Reg.scala 15:16]
  reg  _T_1497; // @[Reg.scala 15:16]
  reg  _T_1498; // @[Reg.scala 15:16]
  reg  _T_1499; // @[Reg.scala 15:16]
  reg  _T_1500; // @[Reg.scala 15:16]
  reg  _T_1501; // @[Reg.scala 15:16]
  reg  _T_1502; // @[Reg.scala 15:16]
  reg  _T_1503; // @[Reg.scala 15:16]
  reg  _T_1504; // @[Reg.scala 15:16]
  reg  _T_1505; // @[Reg.scala 15:16]
  reg  _T_1506; // @[Reg.scala 15:16]
  reg  _T_1507; // @[Reg.scala 15:16]
  reg  _T_1508; // @[Reg.scala 15:16]
  reg  _T_1509; // @[Reg.scala 15:16]
  reg  _T_1510; // @[Reg.scala 15:16]
  reg  _T_1511; // @[Reg.scala 15:16]
  reg  _T_1512; // @[Reg.scala 15:16]
  reg  _T_1513; // @[Reg.scala 15:16]
  reg  _T_1514; // @[Reg.scala 15:16]
  reg  _T_1515; // @[Reg.scala 15:16]
  reg  _T_1516; // @[Reg.scala 15:16]
  reg  _T_1517; // @[Reg.scala 15:16]
  reg  _T_1518; // @[Reg.scala 15:16]
  reg  _T_1519; // @[Reg.scala 15:16]
  reg  _T_1520; // @[Reg.scala 15:16]
  reg  _T_1521; // @[Reg.scala 15:16]
  reg  _T_1522; // @[Reg.scala 15:16]
  reg  _T_1523; // @[Reg.scala 15:16]
  reg  _T_1524; // @[Reg.scala 15:16]
  reg  _T_1525; // @[Reg.scala 15:16]
  reg  _T_1526; // @[Reg.scala 15:16]
  reg  _T_1527; // @[Reg.scala 15:16]
  reg  _T_1528; // @[Reg.scala 15:16]
  reg  _T_1529; // @[Reg.scala 15:16]
  reg  _T_1530; // @[Reg.scala 15:16]
  reg  _T_1531; // @[Reg.scala 15:16]
  reg  _T_1532; // @[Reg.scala 15:16]
  reg  _T_1533; // @[Reg.scala 15:16]
  reg  _T_1534; // @[Reg.scala 15:16]
  reg  _T_1535; // @[Reg.scala 15:16]
  reg  _T_1536; // @[Reg.scala 15:16]
  reg  _T_1537; // @[Reg.scala 15:16]
  reg  _T_1538; // @[Reg.scala 15:16]
  reg  _T_1539; // @[Reg.scala 15:16]
  reg  _T_1540; // @[Reg.scala 15:16]
  reg  _T_1541; // @[Reg.scala 15:16]
  reg  _T_1542; // @[Reg.scala 15:16]
  reg  _T_1543; // @[Reg.scala 15:16]
  reg  _T_1544; // @[Reg.scala 15:16]
  reg  _T_1545; // @[Reg.scala 15:16]
  reg  _T_1546; // @[Reg.scala 15:16]
  reg  _T_1547; // @[Reg.scala 15:16]
  reg  _T_1548; // @[Reg.scala 15:16]
  reg  _T_1549; // @[Reg.scala 15:16]
  reg  _T_1550; // @[Reg.scala 15:16]
  reg  _T_1551; // @[Reg.scala 15:16]
  reg  _T_1552; // @[Reg.scala 15:16]
  reg  _T_1553; // @[Reg.scala 15:16]
  reg  _T_1554; // @[Reg.scala 15:16]
  reg  _T_1555; // @[Reg.scala 15:16]
  reg  _T_1556; // @[Reg.scala 15:16]
  reg  _T_1557; // @[Reg.scala 15:16]
  reg  _T_1558; // @[Reg.scala 15:16]
  reg  _T_1559; // @[Reg.scala 15:16]
  reg  _T_1560; // @[Reg.scala 15:16]
  reg  _T_1561; // @[Reg.scala 15:16]
  reg  _T_1562; // @[Reg.scala 15:16]
  reg  _T_1563; // @[Reg.scala 15:16]
  reg  _T_1564; // @[Reg.scala 15:16]
  reg  _T_1565; // @[Reg.scala 15:16]
  reg  _T_1566; // @[Reg.scala 15:16]
  reg  _T_1567; // @[Reg.scala 15:16]
  reg  _T_1568; // @[Reg.scala 15:16]
  reg  _T_1569; // @[Reg.scala 15:16]
  reg  _T_1570; // @[Reg.scala 15:16]
  reg  _T_1571; // @[Reg.scala 15:16]
  reg  _T_1572; // @[Reg.scala 15:16]
  reg  _T_1573; // @[Reg.scala 15:16]
  reg  _T_1574; // @[Reg.scala 15:16]
  reg  _T_1575; // @[Reg.scala 15:16]
  reg  _T_1576; // @[Reg.scala 15:16]
  reg  _T_1577; // @[Reg.scala 15:16]
  reg  _T_1578; // @[Reg.scala 15:16]
  reg  _T_1579; // @[Reg.scala 15:16]
  reg  _T_1580; // @[Reg.scala 15:16]
  reg  _T_1581; // @[Reg.scala 15:16]
  reg  _T_1582; // @[Reg.scala 15:16]
  reg  _T_1583; // @[Reg.scala 15:16]
  reg  _T_1584; // @[Reg.scala 15:16]
  reg  _T_1585; // @[Reg.scala 15:16]
  reg  _T_1586; // @[Reg.scala 15:16]
  reg  _T_1587; // @[Reg.scala 15:16]
  reg  _T_1588; // @[Reg.scala 15:16]
  reg  _T_1589; // @[Reg.scala 15:16]
  reg  _T_1590; // @[Reg.scala 15:16]
  reg  _T_1591; // @[Reg.scala 15:16]
  reg  _T_1592; // @[Reg.scala 15:16]
  reg  _T_1593; // @[Reg.scala 15:16]
  reg  _T_1594; // @[Reg.scala 15:16]
  reg  _T_1595; // @[Reg.scala 15:16]
  reg  _T_1596; // @[Reg.scala 15:16]
  reg  _T_1597; // @[Reg.scala 15:16]
  reg  _T_1598; // @[Reg.scala 15:16]
  reg  _T_1599; // @[Reg.scala 15:16]
  reg  _T_1600; // @[Reg.scala 15:16]
  reg  _T_1601; // @[Reg.scala 15:16]
  reg  _T_1602; // @[Reg.scala 15:16]
  reg  _T_1603; // @[Reg.scala 15:16]
  reg  _T_1604; // @[Reg.scala 15:16]
  reg  _T_1605; // @[Reg.scala 15:16]
  reg  _T_1606; // @[Reg.scala 15:16]
  reg  _T_1607; // @[Reg.scala 15:16]
  reg  _T_1608; // @[Reg.scala 15:16]
  reg  _T_1609; // @[Reg.scala 15:16]
  reg  _T_1610; // @[Reg.scala 15:16]
  reg  _T_1611; // @[Reg.scala 15:16]
  reg  _T_1612; // @[Reg.scala 15:16]
  reg  _T_1613; // @[Reg.scala 15:16]
  reg  _T_1614; // @[Reg.scala 15:16]
  reg  _T_1615; // @[Reg.scala 15:16]
  reg  _T_1616; // @[Reg.scala 15:16]
  reg  _T_1617; // @[Reg.scala 15:16]
  reg  _T_1618; // @[Reg.scala 15:16]
  reg  _T_1619; // @[Reg.scala 15:16]
  reg  _T_1620; // @[Reg.scala 15:16]
  reg  _T_1621; // @[Reg.scala 15:16]
  reg  _T_1622; // @[Reg.scala 15:16]
  reg  _T_1623; // @[Reg.scala 15:16]
  reg  _T_1624; // @[Reg.scala 15:16]
  reg  _T_1625; // @[Reg.scala 15:16]
  reg  _T_1626; // @[Reg.scala 15:16]
  reg  _T_1627; // @[Reg.scala 15:16]
  reg  _T_1628; // @[Reg.scala 15:16]
  reg  _T_1629; // @[Reg.scala 15:16]
  reg  _T_1630; // @[Reg.scala 15:16]
  reg  _T_1631; // @[Reg.scala 15:16]
  reg  _T_1632; // @[Reg.scala 15:16]
  reg  _T_1633; // @[Reg.scala 15:16]
  reg  _T_1634; // @[Reg.scala 15:16]
  reg  _T_1635; // @[Reg.scala 15:16]
  reg  _T_1636; // @[Reg.scala 15:16]
  reg  _T_1637; // @[Reg.scala 15:16]
  reg  _T_1638; // @[Reg.scala 15:16]
  reg  _T_1639; // @[Reg.scala 15:16]
  reg  _T_1640; // @[Reg.scala 15:16]
  reg  _T_1641; // @[Reg.scala 15:16]
  reg  _T_1642; // @[Reg.scala 15:16]
  reg  _T_1643; // @[Reg.scala 15:16]
  reg  _T_1644; // @[Reg.scala 15:16]
  reg  _T_1645; // @[Reg.scala 15:16]
  reg  _T_1646; // @[Reg.scala 15:16]
  reg  _T_1647; // @[Reg.scala 15:16]
  reg  _T_1648; // @[Reg.scala 15:16]
  reg  _T_1649; // @[Reg.scala 15:16]
  reg  _T_1650; // @[Reg.scala 15:16]
  reg  _T_1651; // @[Reg.scala 15:16]
  reg  _T_1652; // @[Reg.scala 15:16]
  reg  _T_1653; // @[Reg.scala 15:16]
  reg  _T_1654; // @[Reg.scala 15:16]
  reg  _T_1655; // @[Reg.scala 15:16]
  reg  _T_1656; // @[Reg.scala 15:16]
  reg  _T_1657; // @[Reg.scala 15:16]
  reg  _T_1658; // @[Reg.scala 15:16]
  reg  _T_1659; // @[Reg.scala 15:16]
  reg  _T_1660; // @[Reg.scala 15:16]
  reg  _T_1661; // @[Reg.scala 15:16]
  reg  _T_1662; // @[Reg.scala 15:16]
  reg  _T_1663; // @[Reg.scala 15:16]
  reg  _T_1664; // @[Reg.scala 15:16]
  reg  _T_1665; // @[Reg.scala 15:16]
  reg  _T_1666; // @[Reg.scala 15:16]
  reg  _T_1667; // @[Reg.scala 15:16]
  reg  _T_1668; // @[Reg.scala 15:16]
  reg  _T_1669; // @[Reg.scala 15:16]
  reg  _T_1670; // @[Reg.scala 15:16]
  reg  _T_1671; // @[Reg.scala 15:16]
  reg  _T_1672; // @[Reg.scala 15:16]
  reg  _T_1673; // @[Reg.scala 15:16]
  reg  _T_1674; // @[Reg.scala 15:16]
  reg  _T_1675; // @[Reg.scala 15:16]
  reg  _T_1676; // @[Reg.scala 15:16]
  reg  _T_1677; // @[Reg.scala 15:16]
  reg  _T_1678; // @[Reg.scala 15:16]
  reg  _T_1679; // @[Reg.scala 15:16]
  reg  _T_1680; // @[Reg.scala 15:16]
  reg  _T_1681; // @[Reg.scala 15:16]
  reg  _T_1682; // @[Reg.scala 15:16]
  reg  _T_1683; // @[Reg.scala 15:16]
  reg  _T_1684; // @[Reg.scala 15:16]
  reg  _T_1685; // @[Reg.scala 15:16]
  reg  _T_1686; // @[Reg.scala 15:16]
  reg  _T_1687; // @[Reg.scala 15:16]
  reg  _T_1688; // @[Reg.scala 15:16]
  reg  _T_1689; // @[Reg.scala 15:16]
  reg  _T_1690; // @[Reg.scala 15:16]
  reg  _T_1691; // @[Reg.scala 15:16]
  reg  _T_1692; // @[Reg.scala 15:16]
  reg  _T_1693; // @[Reg.scala 15:16]
  reg  _T_1694; // @[Reg.scala 15:16]
  reg  _T_1695; // @[Reg.scala 15:16]
  reg  _T_1696; // @[Reg.scala 15:16]
  reg  _T_1697; // @[Reg.scala 15:16]
  reg  _T_1698; // @[Reg.scala 15:16]
  reg  _T_1699; // @[Reg.scala 15:16]
  reg  _T_1700; // @[Reg.scala 15:16]
  reg  _T_1701; // @[Reg.scala 15:16]
  reg  _T_1702; // @[Reg.scala 15:16]
  reg  _T_1703; // @[Reg.scala 15:16]
  reg  _T_1704; // @[Reg.scala 15:16]
  reg  _T_1705; // @[Reg.scala 15:16]
  reg  _T_1706; // @[Reg.scala 15:16]
  reg  _T_1707; // @[Reg.scala 15:16]
  reg  _T_1708; // @[Reg.scala 15:16]
  reg  _T_1709; // @[Reg.scala 15:16]
  reg  _T_1710; // @[Reg.scala 15:16]
  reg  _T_1711; // @[Reg.scala 15:16]
  reg  _T_1712; // @[Reg.scala 15:16]
  reg  _T_1713; // @[Reg.scala 15:16]
  reg  _T_1714; // @[Reg.scala 15:16]
  reg  _T_1715; // @[Reg.scala 15:16]
  reg  _T_1716; // @[Reg.scala 15:16]
  reg  _T_1717; // @[Reg.scala 15:16]
  reg  _T_1718; // @[Reg.scala 15:16]
  reg  _T_1719; // @[Reg.scala 15:16]
  reg  _T_1720; // @[Reg.scala 15:16]
  reg  _T_1721; // @[Reg.scala 15:16]
  reg  _T_1722; // @[Reg.scala 15:16]
  reg  _T_1723; // @[Reg.scala 15:16]
  reg  _T_1724; // @[Reg.scala 15:16]
  reg  _T_1725; // @[Reg.scala 15:16]
  reg  _T_1726; // @[Reg.scala 15:16]
  reg  _T_1727; // @[Reg.scala 15:16]
  reg  _T_1728; // @[Reg.scala 15:16]
  reg  _T_1729; // @[Reg.scala 15:16]
  reg  _T_1730; // @[Reg.scala 15:16]
  reg  _T_1731; // @[Reg.scala 15:16]
  reg  _T_1732; // @[Reg.scala 15:16]
  reg  _T_1733; // @[Reg.scala 15:16]
  reg  _T_1734; // @[Reg.scala 15:16]
  reg  _T_1735; // @[Reg.scala 15:16]
  reg  _T_1736; // @[Reg.scala 15:16]
  reg  _T_1737; // @[Reg.scala 15:16]
  reg  _T_1738; // @[Reg.scala 15:16]
  reg  _T_1739; // @[Reg.scala 15:16]
  reg  _T_1740; // @[Reg.scala 15:16]
  reg  _T_1741; // @[Reg.scala 15:16]
  reg  _T_1742; // @[Reg.scala 15:16]
  reg  _T_1743; // @[Reg.scala 15:16]
  reg  _T_1744; // @[Reg.scala 15:16]
  reg  _T_1745; // @[Reg.scala 15:16]
  reg  _T_1746; // @[Reg.scala 15:16]
  reg  _T_1747; // @[Reg.scala 15:16]
  reg  _T_1748; // @[Reg.scala 15:16]
  reg  _T_1749; // @[Reg.scala 15:16]
  reg  _T_1750; // @[Reg.scala 15:16]
  reg  _T_1751; // @[Reg.scala 15:16]
  reg  _T_1752; // @[Reg.scala 15:16]
  reg  _T_1753; // @[Reg.scala 15:16]
  reg  _T_1754; // @[Reg.scala 15:16]
  reg  _T_1755; // @[Reg.scala 15:16]
  reg  _T_1756; // @[Reg.scala 15:16]
  reg  _T_1757; // @[Reg.scala 15:16]
  reg  _T_1758; // @[Reg.scala 15:16]
  reg  _T_1759; // @[Reg.scala 15:16]
  reg  _T_1760; // @[Reg.scala 15:16]
  reg  _T_1761; // @[Reg.scala 15:16]
  reg  _T_1762; // @[Reg.scala 15:16]
  reg  _T_1763; // @[Reg.scala 15:16]
  reg  _T_1764; // @[Reg.scala 15:16]
  reg  _T_1765; // @[Reg.scala 15:16]
  reg  _T_1766; // @[Reg.scala 15:16]
  reg  _T_1767; // @[Reg.scala 15:16]
  reg  _T_1768; // @[Reg.scala 15:16]
  reg  _T_1769; // @[Reg.scala 15:16]
  reg  _T_1770; // @[Reg.scala 15:16]
  reg  _T_1771; // @[Reg.scala 15:16]
  reg  _T_1772; // @[Reg.scala 15:16]
  reg  _T_1773; // @[Reg.scala 15:16]
  reg  _T_1774; // @[Reg.scala 15:16]
  reg  _T_1775; // @[Reg.scala 15:16]
  reg  _T_1776; // @[Reg.scala 15:16]
  reg  _T_1777; // @[Reg.scala 15:16]
  reg  _T_1778; // @[Reg.scala 15:16]
  reg  _T_1779; // @[Reg.scala 15:16]
  reg  _T_1780; // @[Reg.scala 15:16]
  reg  _T_1781; // @[Reg.scala 15:16]
  reg  _T_1782; // @[Reg.scala 15:16]
  reg  _T_1783; // @[Reg.scala 15:16]
  reg  _T_1784; // @[Reg.scala 15:16]
  reg  _T_1785; // @[Reg.scala 15:16]
  reg  _T_1786; // @[Reg.scala 15:16]
  reg  _T_1787; // @[Reg.scala 15:16]
  reg  _T_1788; // @[Reg.scala 15:16]
  reg  _T_1789; // @[Reg.scala 15:16]
  reg  _T_1790; // @[Reg.scala 15:16]
  reg  _T_1791; // @[Reg.scala 15:16]
  reg  _T_1792; // @[Reg.scala 15:16]
  reg  _T_1793; // @[Reg.scala 15:16]
  reg  _T_1794; // @[Reg.scala 15:16]
  reg  _T_1795; // @[Reg.scala 15:16]
  reg  _T_1796; // @[Reg.scala 15:16]
  reg  _T_1797; // @[Reg.scala 15:16]
  reg  _T_1798; // @[Reg.scala 15:16]
  reg  _T_1799; // @[Reg.scala 15:16]
  reg  _T_1800; // @[Reg.scala 15:16]
  reg  _T_1801; // @[Reg.scala 15:16]
  reg  _T_1802; // @[Reg.scala 15:16]
  reg  _T_1803; // @[Reg.scala 15:16]
  reg  _T_1804; // @[Reg.scala 15:16]
  reg  _T_1805; // @[Reg.scala 15:16]
  reg  _T_1806; // @[Reg.scala 15:16]
  reg  _T_1807; // @[Reg.scala 15:16]
  reg  _T_1808; // @[Reg.scala 15:16]
  reg  _T_1809; // @[Reg.scala 15:16]
  reg  _T_1810; // @[Reg.scala 15:16]
  reg  _T_1811; // @[Reg.scala 15:16]
  reg  _T_1812; // @[Reg.scala 15:16]
  reg  _T_1813; // @[Reg.scala 15:16]
  reg  _T_1814; // @[Reg.scala 15:16]
  reg  _T_1815; // @[Reg.scala 15:16]
  reg  _T_1816; // @[Reg.scala 15:16]
  reg  _T_1817; // @[Reg.scala 15:16]
  reg  _T_1818; // @[Reg.scala 15:16]
  reg  _T_1819; // @[Reg.scala 15:16]
  reg  _T_1820; // @[Reg.scala 15:16]
  reg  _T_1821; // @[Reg.scala 15:16]
  reg  _T_1822; // @[Reg.scala 15:16]
  reg  _T_1823; // @[Reg.scala 15:16]
  reg  _T_1824; // @[Reg.scala 15:16]
  reg  _T_1825; // @[Reg.scala 15:16]
  reg  _T_1826; // @[Reg.scala 15:16]
  reg  _T_1827; // @[Reg.scala 15:16]
  reg  _T_1828; // @[Reg.scala 15:16]
  reg  _T_1829; // @[Reg.scala 15:16]
  reg  _T_1830; // @[Reg.scala 15:16]
  reg  _T_1831; // @[Reg.scala 15:16]
  reg  _T_1832; // @[Reg.scala 15:16]
  reg  _T_1833; // @[Reg.scala 15:16]
  reg  _T_1834; // @[Reg.scala 15:16]
  reg  _T_1835; // @[Reg.scala 15:16]
  reg  _T_1836; // @[Reg.scala 15:16]
  reg  _T_1837; // @[Reg.scala 15:16]
  reg  _T_1838; // @[Reg.scala 15:16]
  reg  _T_1839; // @[Reg.scala 15:16]
  reg  _T_1840; // @[Reg.scala 15:16]
  reg  _T_1841; // @[Reg.scala 15:16]
  reg  _T_1842; // @[Reg.scala 15:16]
  reg  _T_1843; // @[Reg.scala 15:16]
  reg  _T_1844; // @[Reg.scala 15:16]
  reg  _T_1845; // @[Reg.scala 15:16]
  reg  _T_1846; // @[Reg.scala 15:16]
  reg  _T_1847; // @[Reg.scala 15:16]
  reg  _T_1848; // @[Reg.scala 15:16]
  reg  _T_1849; // @[Reg.scala 15:16]
  reg  _T_1850; // @[Reg.scala 15:16]
  reg  _T_1851; // @[Reg.scala 15:16]
  reg  _T_1852; // @[Reg.scala 15:16]
  reg  _T_1853; // @[Reg.scala 15:16]
  reg  _T_1854; // @[Reg.scala 15:16]
  reg  _T_1855; // @[Reg.scala 15:16]
  reg  _T_1856; // @[Reg.scala 15:16]
  reg  _T_1857; // @[Reg.scala 15:16]
  reg  _T_1858; // @[Reg.scala 15:16]
  reg  _T_1859; // @[Reg.scala 15:16]
  reg  _T_1860; // @[Reg.scala 15:16]
  reg  _T_1861; // @[Reg.scala 15:16]
  reg  _T_1862; // @[Reg.scala 15:16]
  reg  _T_1863; // @[Reg.scala 15:16]
  reg  _T_1864; // @[Reg.scala 15:16]
  reg  _T_1865; // @[Reg.scala 15:16]
  reg  _T_1866; // @[Reg.scala 15:16]
  reg  _T_1867; // @[Reg.scala 15:16]
  reg  _T_1868; // @[Reg.scala 15:16]
  reg  _T_1869; // @[Reg.scala 15:16]
  reg  _T_1870; // @[Reg.scala 15:16]
  reg  _T_1871; // @[Reg.scala 15:16]
  reg  _T_1872; // @[Reg.scala 15:16]
  reg  _T_1873; // @[Reg.scala 15:16]
  reg  _T_1874; // @[Reg.scala 15:16]
  reg  _T_1875; // @[Reg.scala 15:16]
  reg  _T_1876; // @[Reg.scala 15:16]
  reg  _T_1877; // @[Reg.scala 15:16]
  reg  _T_1878; // @[Reg.scala 15:16]
  reg  _T_1879; // @[Reg.scala 15:16]
  reg  _T_1880; // @[Reg.scala 15:16]
  reg  _T_1881; // @[Reg.scala 15:16]
  reg  _T_1882; // @[Reg.scala 15:16]
  reg  _T_1883; // @[Reg.scala 15:16]
  reg  _T_1884; // @[Reg.scala 15:16]
  reg  _T_1885; // @[Reg.scala 15:16]
  reg  _T_1886; // @[Reg.scala 15:16]
  reg  _T_1887; // @[Reg.scala 15:16]
  reg  _T_1888; // @[Reg.scala 15:16]
  reg  _T_1889; // @[Reg.scala 15:16]
  reg  _T_1890; // @[Reg.scala 15:16]
  reg  _T_1891; // @[Reg.scala 15:16]
  reg  _T_1892; // @[Reg.scala 15:16]
  reg  _T_1893; // @[Reg.scala 15:16]
  reg  _T_1894; // @[Reg.scala 15:16]
  reg  _T_1895; // @[Reg.scala 15:16]
  reg  _T_1896; // @[Reg.scala 15:16]
  reg  _T_1897; // @[Reg.scala 15:16]
  reg  _T_1898; // @[Reg.scala 15:16]
  reg  _T_1899; // @[Reg.scala 15:16]
  reg  _T_1900; // @[Reg.scala 15:16]
  reg  _T_1901; // @[Reg.scala 15:16]
  reg  _T_1902; // @[Reg.scala 15:16]
  reg  _T_1903; // @[Reg.scala 15:16]
  reg  _T_1904; // @[Reg.scala 15:16]
  reg  _T_1905; // @[Reg.scala 15:16]
  reg  _T_1906; // @[Reg.scala 15:16]
  reg  _T_1907; // @[Reg.scala 15:16]
  reg  _T_1908; // @[Reg.scala 15:16]
  reg  _T_1909; // @[Reg.scala 15:16]
  reg  _T_1910; // @[Reg.scala 15:16]
  reg  _T_1911; // @[Reg.scala 15:16]
  reg  _T_1912; // @[Reg.scala 15:16]
  reg  _T_1913; // @[Reg.scala 15:16]
  reg  _T_1914; // @[Reg.scala 15:16]
  reg  _T_1915; // @[Reg.scala 15:16]
  reg  _T_1916; // @[Reg.scala 15:16]
  reg  _T_1917; // @[Reg.scala 15:16]
  reg  _T_1918; // @[Reg.scala 15:16]
  reg  _T_1919; // @[Reg.scala 15:16]
  reg  _T_1920; // @[Reg.scala 15:16]
  reg  _T_1921; // @[Reg.scala 15:16]
  reg  _T_1922; // @[Reg.scala 15:16]
  reg  _T_1923; // @[Reg.scala 15:16]
  reg  _T_1924; // @[Reg.scala 15:16]
  reg  _T_1925; // @[Reg.scala 15:16]
  reg  _T_1926; // @[Reg.scala 15:16]
  reg  _T_1927; // @[Reg.scala 15:16]
  reg  _T_1928; // @[Reg.scala 15:16]
  reg  _T_1929; // @[Reg.scala 15:16]
  reg  _T_1930; // @[Reg.scala 15:16]
  reg  _T_1931; // @[Reg.scala 15:16]
  reg  _T_1932; // @[Reg.scala 15:16]
  reg  _T_1933; // @[Reg.scala 15:16]
  reg  _T_1934; // @[Reg.scala 15:16]
  reg  _T_1935; // @[Reg.scala 15:16]
  reg  _T_1936; // @[Reg.scala 15:16]
  reg  _T_1937; // @[Reg.scala 15:16]
  reg  _T_1938; // @[Reg.scala 15:16]
  reg  _T_1939; // @[Reg.scala 15:16]
  reg  _T_1940; // @[Reg.scala 15:16]
  reg  _T_1941; // @[Reg.scala 15:16]
  reg  _T_1942; // @[Reg.scala 15:16]
  reg  _T_1943; // @[Reg.scala 15:16]
  reg  _T_1944; // @[Reg.scala 15:16]
  reg  _T_1945; // @[Reg.scala 15:16]
  reg  _T_1946; // @[Reg.scala 15:16]
  reg  _T_1947; // @[Reg.scala 15:16]
  reg  _T_1948; // @[Reg.scala 15:16]
  reg  _T_1949; // @[Reg.scala 15:16]
  reg  _T_1950; // @[Reg.scala 15:16]
  reg  _T_1951; // @[Reg.scala 15:16]
  reg  _T_1952; // @[Reg.scala 15:16]
  reg  _T_1953; // @[Reg.scala 15:16]
  reg  _T_1954; // @[Reg.scala 15:16]
  reg  _T_1955; // @[Reg.scala 15:16]
  reg  _T_1956; // @[Reg.scala 15:16]
  reg  _T_1957; // @[Reg.scala 15:16]
  reg  _T_1958; // @[Reg.scala 15:16]
  reg  _T_1959; // @[Reg.scala 15:16]
  reg  _T_1960; // @[Reg.scala 15:16]
  reg  _T_1961; // @[Reg.scala 15:16]
  reg  _T_1962; // @[Reg.scala 15:16]
  reg  _T_1963; // @[Reg.scala 15:16]
  reg  _T_1964; // @[Reg.scala 15:16]
  reg  _T_1965; // @[Reg.scala 15:16]
  reg  _T_1966; // @[Reg.scala 15:16]
  reg  _T_1967; // @[Reg.scala 15:16]
  reg  _T_1968; // @[Reg.scala 15:16]
  reg  _T_1969; // @[Reg.scala 15:16]
  reg  _T_1970; // @[Reg.scala 15:16]
  reg  _T_1971; // @[Reg.scala 15:16]
  reg  _T_1972; // @[Reg.scala 15:16]
  reg  _T_1973; // @[Reg.scala 15:16]
  reg  _T_1974; // @[Reg.scala 15:16]
  reg  _T_1975; // @[Reg.scala 15:16]
  reg  _T_1976; // @[Reg.scala 15:16]
  reg  _T_1977; // @[Reg.scala 15:16]
  reg  _T_1978; // @[Reg.scala 15:16]
  reg  _T_1979; // @[Reg.scala 15:16]
  reg  _T_1980; // @[Reg.scala 15:16]
  reg  _T_1981; // @[Reg.scala 15:16]
  reg  _T_1982; // @[Reg.scala 15:16]
  reg  _T_1983; // @[Reg.scala 15:16]
  reg  _T_1984; // @[Reg.scala 15:16]
  reg  _T_1985; // @[Reg.scala 15:16]
  reg  _T_1986; // @[Reg.scala 15:16]
  reg  _T_1987; // @[Reg.scala 15:16]
  reg  _T_1988; // @[Reg.scala 15:16]
  reg  _T_1989; // @[Reg.scala 15:16]
  reg  _T_1990; // @[Reg.scala 15:16]
  reg  _T_1991; // @[Reg.scala 15:16]
  reg  _T_1992; // @[Reg.scala 15:16]
  reg  _T_1993; // @[Reg.scala 15:16]
  reg  _T_1994; // @[Reg.scala 15:16]
  reg  _T_1995; // @[Reg.scala 15:16]
  reg  _T_1996; // @[Reg.scala 15:16]
  reg  _T_1997; // @[Reg.scala 15:16]
  reg  _T_1998; // @[Reg.scala 15:16]
  reg  _T_1999; // @[Reg.scala 15:16]
  reg  _T_2000; // @[Reg.scala 15:16]
  reg  _T_2001; // @[Reg.scala 15:16]
  reg  _T_2002; // @[Reg.scala 15:16]
  reg  _T_2003; // @[Reg.scala 15:16]
  reg  _T_2004; // @[Reg.scala 15:16]
  reg  _T_2005; // @[Reg.scala 15:16]
  reg  _T_2006; // @[Reg.scala 15:16]
  reg  _T_2007; // @[Reg.scala 15:16]
  reg  _T_2008; // @[Reg.scala 15:16]
  reg  _T_2009; // @[Reg.scala 15:16]
  reg  _T_2010; // @[Reg.scala 15:16]
  reg  _T_2011; // @[Reg.scala 15:16]
  reg  _T_2012; // @[Reg.scala 15:16]
  reg  _T_2013; // @[Reg.scala 15:16]
  reg  _T_2014; // @[Reg.scala 15:16]
  reg  _T_2015; // @[Reg.scala 15:16]
  reg  _T_2016; // @[Reg.scala 15:16]
  reg  _T_2017; // @[Reg.scala 15:16]
  reg  _T_2018; // @[Reg.scala 15:16]
  reg  _T_2019; // @[Reg.scala 15:16]
  reg  _T_2020; // @[Reg.scala 15:16]
  reg  _T_2021; // @[Reg.scala 15:16]
  reg  _T_2022; // @[Reg.scala 15:16]
  reg  _T_2023; // @[Reg.scala 15:16]
  reg  _T_2024; // @[Reg.scala 15:16]
  reg  _T_2025; // @[Reg.scala 15:16]
  reg  _T_2026; // @[Reg.scala 15:16]
  reg  _T_2027; // @[Reg.scala 15:16]
  reg  _T_2028; // @[Reg.scala 15:16]
  reg  _T_2029; // @[Reg.scala 15:16]
  reg  _T_2030; // @[Reg.scala 15:16]
  reg  _T_2031; // @[Reg.scala 15:16]
  reg  _T_2032; // @[Reg.scala 15:16]
  reg  _T_2033; // @[Reg.scala 15:16]
  reg  _T_2034; // @[Reg.scala 15:16]
  reg  _T_2035; // @[Reg.scala 15:16]
  reg  _T_2036; // @[Reg.scala 15:16]
  reg  _T_2037; // @[Reg.scala 15:16]
  reg  _T_2038; // @[Reg.scala 15:16]
  reg  _T_2039; // @[Reg.scala 15:16]
  reg  _T_2040; // @[Reg.scala 15:16]
  reg  _T_2041; // @[Reg.scala 15:16]
  reg  _T_2042; // @[Reg.scala 15:16]
  reg  _T_2043; // @[Reg.scala 15:16]
  reg  _T_2044; // @[Reg.scala 15:16]
  reg  _T_2045; // @[Reg.scala 15:16]
  reg  _T_2046; // @[Reg.scala 15:16]
  reg  _T_2047; // @[Reg.scala 15:16]
  reg  _T_2048; // @[Reg.scala 15:16]
  reg  _T_2049; // @[Reg.scala 15:16]
  reg  _T_2050; // @[Reg.scala 15:16]
  reg  _T_2051; // @[Reg.scala 15:16]
  reg  _T_2052; // @[Reg.scala 15:16]
  reg  _T_2053; // @[Reg.scala 15:16]
  reg  _T_2054; // @[Reg.scala 15:16]
  reg  _T_2055; // @[Reg.scala 15:16]
  reg  _T_2056; // @[Reg.scala 15:16]
  reg  _T_2057; // @[Reg.scala 15:16]
  reg  _T_2058; // @[Reg.scala 15:16]
  reg  _T_2059; // @[Reg.scala 15:16]
  reg  _T_2060; // @[Reg.scala 15:16]
  reg  _T_2061; // @[Reg.scala 15:16]
  reg  _T_2062; // @[Reg.scala 15:16]
  reg  _T_2063; // @[Reg.scala 15:16]
  reg  _T_2064; // @[Reg.scala 15:16]
  reg  _T_2065; // @[Reg.scala 15:16]
  reg  _T_2066; // @[Reg.scala 15:16]
  reg  _T_2067; // @[Reg.scala 15:16]
  reg  _T_2068; // @[Reg.scala 15:16]
  reg  _T_2069; // @[Reg.scala 15:16]
  reg  _T_2070; // @[Reg.scala 15:16]
  reg  _T_2071; // @[Reg.scala 15:16]
  reg  _T_2072; // @[Reg.scala 15:16]
  reg  _T_2073; // @[Reg.scala 15:16]
  reg  _T_2074; // @[Reg.scala 15:16]
  reg  _T_2075; // @[Reg.scala 15:16]
  reg  _T_2076; // @[Reg.scala 15:16]
  reg  _T_2077; // @[Reg.scala 15:16]
  reg  _T_2078; // @[Reg.scala 15:16]
  reg  _T_2079; // @[Reg.scala 15:16]
  reg  _T_2080; // @[Reg.scala 15:16]
  reg  _T_2081; // @[Reg.scala 15:16]
  reg  _T_2082; // @[Reg.scala 15:16]
  reg  _T_2083; // @[Reg.scala 15:16]
  reg  _T_2084; // @[Reg.scala 15:16]
  reg  _T_2085; // @[Reg.scala 15:16]
  reg  _T_2086; // @[Reg.scala 15:16]
  reg  _T_2087; // @[Reg.scala 15:16]
  reg  _T_2088; // @[Reg.scala 15:16]
  reg  _T_2089; // @[Reg.scala 15:16]
  reg  _T_2090; // @[Reg.scala 15:16]
  reg  _T_2091; // @[Reg.scala 15:16]
  reg  _T_2092; // @[Reg.scala 15:16]
  reg  _T_2093; // @[Reg.scala 15:16]
  reg  _T_2094; // @[Reg.scala 15:16]
  reg  _T_2095; // @[Reg.scala 15:16]
  reg  _T_2096; // @[Reg.scala 15:16]
  reg  _T_2097; // @[Reg.scala 15:16]
  reg  _T_2098; // @[Reg.scala 15:16]
  reg  _T_2099; // @[Reg.scala 15:16]
  reg  _T_2100; // @[Reg.scala 15:16]
  reg  _T_2101; // @[Reg.scala 15:16]
  reg  _T_2102; // @[Reg.scala 15:16]
  reg  _T_2103; // @[Reg.scala 15:16]
  reg  _T_2104; // @[Reg.scala 15:16]
  reg  _T_2105; // @[Reg.scala 15:16]
  reg  _T_2106; // @[Reg.scala 15:16]
  reg  _T_2107; // @[Reg.scala 15:16]
  reg  _T_2108; // @[Reg.scala 15:16]
  reg  _T_2109; // @[Reg.scala 15:16]
  reg  _T_2110; // @[Reg.scala 15:16]
  reg  _T_2111; // @[Reg.scala 15:16]
  reg  _T_2112; // @[Reg.scala 15:16]
  reg  _T_2113; // @[Reg.scala 15:16]
  reg  _T_2114; // @[Reg.scala 15:16]
  reg  _T_2115; // @[Reg.scala 15:16]
  reg  _T_2116; // @[Reg.scala 15:16]
  reg  _T_2117; // @[Reg.scala 15:16]
  reg  _T_2118; // @[Reg.scala 15:16]
  reg  _T_2119; // @[Reg.scala 15:16]
  reg  _T_2120; // @[Reg.scala 15:16]
  reg  _T_2121; // @[Reg.scala 15:16]
  reg  _T_2122; // @[Reg.scala 15:16]
  reg  _T_2123; // @[Reg.scala 15:16]
  reg  _T_2124; // @[Reg.scala 15:16]
  reg  _T_2125; // @[Reg.scala 15:16]
  reg  _T_2126; // @[Reg.scala 15:16]
  reg  _T_2127; // @[Reg.scala 15:16]
  reg  _T_2128; // @[Reg.scala 15:16]
  reg  _T_2129; // @[Reg.scala 15:16]
  reg  _T_2130; // @[Reg.scala 15:16]
  reg  _T_2131; // @[Reg.scala 15:16]
  reg  _T_2132; // @[Reg.scala 15:16]
  reg  _T_2133; // @[Reg.scala 15:16]
  reg  _T_2134; // @[Reg.scala 15:16]
  reg  _T_2135; // @[Reg.scala 15:16]
  reg  _T_2136; // @[Reg.scala 15:16]
  reg  _T_2137; // @[Reg.scala 15:16]
  reg  _T_2138; // @[Reg.scala 15:16]
  reg  _T_2139; // @[Reg.scala 15:16]
  reg  _T_2140; // @[Reg.scala 15:16]
  reg  _T_2141; // @[Reg.scala 15:16]
  reg  _T_2142; // @[Reg.scala 15:16]
  reg  _T_2143; // @[Reg.scala 15:16]
  reg  _T_2144; // @[Reg.scala 15:16]
  reg  _T_2145; // @[Reg.scala 15:16]
  reg  _T_2146; // @[Reg.scala 15:16]
  reg  _T_2147; // @[Reg.scala 15:16]
  reg  _T_2148; // @[Reg.scala 15:16]
  reg  _T_2149; // @[Reg.scala 15:16]
  reg  _T_2150; // @[Reg.scala 15:16]
  reg  _T_2151; // @[Reg.scala 15:16]
  reg  _T_2152; // @[Reg.scala 15:16]
  reg  _T_2153; // @[Reg.scala 15:16]
  reg  _T_2154; // @[Reg.scala 15:16]
  reg  _T_2155; // @[Reg.scala 15:16]
  reg  _T_2156; // @[Reg.scala 15:16]
  reg  _T_2157; // @[Reg.scala 15:16]
  reg  _T_2158; // @[Reg.scala 15:16]
  reg  _T_2159; // @[Reg.scala 15:16]
  reg  _T_2160; // @[Reg.scala 15:16]
  reg  _T_2161; // @[Reg.scala 15:16]
  reg  _T_2162; // @[Reg.scala 15:16]
  reg  _T_2163; // @[Reg.scala 15:16]
  reg  _T_2164; // @[Reg.scala 15:16]
  reg  _T_2165; // @[Reg.scala 15:16]
  reg  _T_2166; // @[Reg.scala 15:16]
  reg  _T_2167; // @[Reg.scala 15:16]
  reg  _T_2168; // @[Reg.scala 15:16]
  reg  _T_2169; // @[Reg.scala 15:16]
  reg  _T_2170; // @[Reg.scala 15:16]
  reg  _T_2171; // @[Reg.scala 15:16]
  reg  _T_2172; // @[Reg.scala 15:16]
  reg  _T_2173; // @[Reg.scala 15:16]
  reg  _T_2174; // @[Reg.scala 15:16]
  reg  _T_2175; // @[Reg.scala 15:16]
  reg  _T_2176; // @[Reg.scala 15:16]
  reg  _T_2177; // @[Reg.scala 15:16]
  reg  _T_2178; // @[Reg.scala 15:16]
  reg  _T_2179; // @[Reg.scala 15:16]
  reg  _T_2180; // @[Reg.scala 15:16]
  reg  _T_2181; // @[Reg.scala 15:16]
  reg  _T_2182; // @[Reg.scala 15:16]
  reg  _T_2183; // @[Reg.scala 15:16]
  reg  _T_2184; // @[Reg.scala 15:16]
  reg  _T_2185; // @[Reg.scala 15:16]
  reg  _T_2186; // @[Reg.scala 15:16]
  reg  _T_2187; // @[Reg.scala 15:16]
  reg  _T_2188; // @[Reg.scala 15:16]
  reg  _T_2189; // @[Reg.scala 15:16]
  reg  _T_2190; // @[Reg.scala 15:16]
  reg  _T_2191; // @[Reg.scala 15:16]
  reg  _T_2192; // @[Reg.scala 15:16]
  reg  _T_2193; // @[Reg.scala 15:16]
  reg  _T_2194; // @[Reg.scala 15:16]
  reg  _T_2195; // @[Reg.scala 15:16]
  reg  _T_2196; // @[Reg.scala 15:16]
  reg  _T_2197; // @[Reg.scala 15:16]
  reg  _T_2198; // @[Reg.scala 15:16]
  reg  _T_2199; // @[Reg.scala 15:16]
  reg  _T_2200; // @[Reg.scala 15:16]
  reg  _T_2201; // @[Reg.scala 15:16]
  reg  _T_2202; // @[Reg.scala 15:16]
  reg  _T_2203; // @[Reg.scala 15:16]
  reg  _T_2204; // @[Reg.scala 15:16]
  reg  _T_2205; // @[Reg.scala 15:16]
  reg  _T_2206; // @[Reg.scala 15:16]
  reg  _T_2207; // @[Reg.scala 15:16]
  reg  _T_2208; // @[Reg.scala 15:16]
  reg  _T_2209; // @[Reg.scala 15:16]
  reg  _T_2210; // @[Reg.scala 15:16]
  reg  _T_2211; // @[Reg.scala 15:16]
  reg  _T_2212; // @[Reg.scala 15:16]
  reg  _T_2213; // @[Reg.scala 15:16]
  reg  _T_2214; // @[Reg.scala 15:16]
  reg  _T_2215; // @[Reg.scala 15:16]
  reg  _T_2216; // @[Reg.scala 15:16]
  reg  _T_2217; // @[Reg.scala 15:16]
  reg  _T_2218; // @[Reg.scala 15:16]
  reg  _T_2219; // @[Reg.scala 15:16]
  reg  _T_2220; // @[Reg.scala 15:16]
  reg  _T_2221; // @[Reg.scala 15:16]
  reg  _T_2222; // @[Reg.scala 15:16]
  reg  _T_2223; // @[Reg.scala 15:16]
  reg  _T_2224; // @[Reg.scala 15:16]
  reg  _T_2225; // @[Reg.scala 15:16]
  reg  _T_2226; // @[Reg.scala 15:16]
  reg  _T_2227; // @[Reg.scala 15:16]
  reg  _T_2228; // @[Reg.scala 15:16]
  reg  _T_2229; // @[Reg.scala 15:16]
  reg  _T_2230; // @[Reg.scala 15:16]
  reg  _T_2231; // @[Reg.scala 15:16]
  reg  _T_2232; // @[Reg.scala 15:16]
  reg  _T_2233; // @[Reg.scala 15:16]
  reg  _T_2234; // @[Reg.scala 15:16]
  reg  _T_2235; // @[Reg.scala 15:16]
  reg  _T_2236; // @[Reg.scala 15:16]
  reg  _T_2237; // @[Reg.scala 15:16]
  reg  _T_2238; // @[Reg.scala 15:16]
  reg  _T_2239; // @[Reg.scala 15:16]
  reg  _T_2240; // @[Reg.scala 15:16]
  reg  _T_2241; // @[Reg.scala 15:16]
  reg  _T_2242; // @[Reg.scala 15:16]
  reg  _T_2243; // @[Reg.scala 15:16]
  reg  _T_2244; // @[Reg.scala 15:16]
  reg  _T_2245; // @[Reg.scala 15:16]
  reg  _T_2246; // @[Reg.scala 15:16]
  reg  _T_2247; // @[Reg.scala 15:16]
  reg  _T_2248; // @[Reg.scala 15:16]
  reg  _T_2249; // @[Reg.scala 15:16]
  reg  _T_2250; // @[Reg.scala 15:16]
  reg  _T_2251; // @[Reg.scala 15:16]
  reg  _T_2252; // @[Reg.scala 15:16]
  reg  _T_2253; // @[Reg.scala 15:16]
  reg  _T_2254; // @[Reg.scala 15:16]
  reg  _T_2255; // @[Reg.scala 15:16]
  reg  _T_2256; // @[Reg.scala 15:16]
  reg  _T_2257; // @[Reg.scala 15:16]
  reg  _T_2258; // @[Reg.scala 15:16]
  reg  _T_2259; // @[Reg.scala 15:16]
  reg  _T_2260; // @[Reg.scala 15:16]
  reg  _T_2261; // @[Reg.scala 15:16]
  reg  _T_2262; // @[Reg.scala 15:16]
  reg  _T_2263; // @[Reg.scala 15:16]
  reg  _T_2264; // @[Reg.scala 15:16]
  reg  _T_2265; // @[Reg.scala 15:16]
  reg  _T_2266; // @[Reg.scala 15:16]
  wire  _T_2267 = ~_T_2266; // @[FFT.scala 90:61]
  Butterfly Butterfly ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_io_in1_re),
    .io_in1_im(Butterfly_io_in1_im),
    .io_in2_re(Butterfly_io_in2_re),
    .io_in2_im(Butterfly_io_in2_im),
    .io_wn_re(Butterfly_io_wn_re),
    .io_wn_im(Butterfly_io_wn_im),
    .io_out1_re(Butterfly_io_out1_re),
    .io_out1_im(Butterfly_io_out1_im),
    .io_out2_re(Butterfly_io_out2_re),
    .io_out2_im(Butterfly_io_out2_im)
  );
  Switch Switch ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  Butterfly Butterfly_1 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_1_io_in1_re),
    .io_in1_im(Butterfly_1_io_in1_im),
    .io_in2_re(Butterfly_1_io_in2_re),
    .io_in2_im(Butterfly_1_io_in2_im),
    .io_wn_re(Butterfly_1_io_wn_re),
    .io_wn_im(Butterfly_1_io_wn_im),
    .io_out1_re(Butterfly_1_io_out1_re),
    .io_out1_im(Butterfly_1_io_out1_im),
    .io_out2_re(Butterfly_1_io_out2_re),
    .io_out2_im(Butterfly_1_io_out2_im)
  );
  Switch Switch_1 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  Butterfly Butterfly_2 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_2_io_in1_re),
    .io_in1_im(Butterfly_2_io_in1_im),
    .io_in2_re(Butterfly_2_io_in2_re),
    .io_in2_im(Butterfly_2_io_in2_im),
    .io_wn_re(Butterfly_2_io_wn_re),
    .io_wn_im(Butterfly_2_io_wn_im),
    .io_out1_re(Butterfly_2_io_out1_re),
    .io_out1_im(Butterfly_2_io_out1_im),
    .io_out2_re(Butterfly_2_io_out2_re),
    .io_out2_im(Butterfly_2_io_out2_im)
  );
  Switch Switch_2 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  Butterfly Butterfly_3 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_3_io_in1_re),
    .io_in1_im(Butterfly_3_io_in1_im),
    .io_in2_re(Butterfly_3_io_in2_re),
    .io_in2_im(Butterfly_3_io_in2_im),
    .io_wn_re(Butterfly_3_io_wn_re),
    .io_wn_im(Butterfly_3_io_wn_im),
    .io_out1_re(Butterfly_3_io_out1_re),
    .io_out1_im(Butterfly_3_io_out1_im),
    .io_out2_re(Butterfly_3_io_out2_re),
    .io_out2_im(Butterfly_3_io_out2_im)
  );
  Switch Switch_3 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  Butterfly Butterfly_4 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_4_io_in1_re),
    .io_in1_im(Butterfly_4_io_in1_im),
    .io_in2_re(Butterfly_4_io_in2_re),
    .io_in2_im(Butterfly_4_io_in2_im),
    .io_wn_re(Butterfly_4_io_wn_re),
    .io_wn_im(Butterfly_4_io_wn_im),
    .io_out1_re(Butterfly_4_io_out1_re),
    .io_out1_im(Butterfly_4_io_out1_im),
    .io_out2_re(Butterfly_4_io_out2_re),
    .io_out2_im(Butterfly_4_io_out2_im)
  );
  Switch Switch_4 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  Butterfly Butterfly_5 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_5_io_in1_re),
    .io_in1_im(Butterfly_5_io_in1_im),
    .io_in2_re(Butterfly_5_io_in2_re),
    .io_in2_im(Butterfly_5_io_in2_im),
    .io_wn_re(Butterfly_5_io_wn_re),
    .io_wn_im(Butterfly_5_io_wn_im),
    .io_out1_re(Butterfly_5_io_out1_re),
    .io_out1_im(Butterfly_5_io_out1_im),
    .io_out2_re(Butterfly_5_io_out2_re),
    .io_out2_im(Butterfly_5_io_out2_im)
  );
  Switch Switch_5 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_5_io_in1_re),
    .io_in1_im(Switch_5_io_in1_im),
    .io_in2_re(Switch_5_io_in2_re),
    .io_in2_im(Switch_5_io_in2_im),
    .io_sel(Switch_5_io_sel),
    .io_out1_re(Switch_5_io_out1_re),
    .io_out1_im(Switch_5_io_out1_im),
    .io_out2_re(Switch_5_io_out2_re),
    .io_out2_im(Switch_5_io_out2_im)
  );
  Butterfly Butterfly_6 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_6_io_in1_re),
    .io_in1_im(Butterfly_6_io_in1_im),
    .io_in2_re(Butterfly_6_io_in2_re),
    .io_in2_im(Butterfly_6_io_in2_im),
    .io_wn_re(Butterfly_6_io_wn_re),
    .io_wn_im(Butterfly_6_io_wn_im),
    .io_out1_re(Butterfly_6_io_out1_re),
    .io_out1_im(Butterfly_6_io_out1_im),
    .io_out2_re(Butterfly_6_io_out2_re),
    .io_out2_im(Butterfly_6_io_out2_im)
  );
  Switch Switch_6 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_6_io_in1_re),
    .io_in1_im(Switch_6_io_in1_im),
    .io_in2_re(Switch_6_io_in2_re),
    .io_in2_im(Switch_6_io_in2_im),
    .io_sel(Switch_6_io_sel),
    .io_out1_re(Switch_6_io_out1_re),
    .io_out1_im(Switch_6_io_out1_im),
    .io_out2_re(Switch_6_io_out2_re),
    .io_out2_im(Switch_6_io_out2_im)
  );
  Butterfly Butterfly_7 ( // @[Butterfly.scala 89:22]
    .io_in1_re(Butterfly_7_io_in1_re),
    .io_in1_im(Butterfly_7_io_in1_im),
    .io_in2_re(Butterfly_7_io_in2_re),
    .io_in2_im(Butterfly_7_io_in2_im),
    .io_wn_re(Butterfly_7_io_wn_re),
    .io_wn_im(Butterfly_7_io_wn_im),
    .io_out1_re(Butterfly_7_io_out1_re),
    .io_out1_im(Butterfly_7_io_out1_im),
    .io_out2_re(Butterfly_7_io_out2_re),
    .io_out2_im(Butterfly_7_io_out2_im)
  );
  Switch Switch_7 ( // @[Butterfly.scala 110:22]
    .io_in1_re(Switch_7_io_in1_re),
    .io_in1_im(Switch_7_io_in1_im),
    .io_in2_re(Switch_7_io_in2_re),
    .io_in2_im(Switch_7_io_in2_im),
    .io_sel(Switch_7_io_sel),
    .io_out1_re(Switch_7_io_out1_re),
    .io_out1_im(Switch_7_io_out1_im),
    .io_out2_re(Switch_7_io_out2_re),
    .io_out2_im(Switch_7_io_out2_im)
  );
  ComplexAdd ComplexAdd ( // @[Butterfly.scala 26:22]
    .io_op1_re(ComplexAdd_io_op1_re),
    .io_op1_im(ComplexAdd_io_op1_im),
    .io_op2_re(ComplexAdd_io_op2_re),
    .io_op2_im(ComplexAdd_io_op2_im),
    .io_res_re(ComplexAdd_io_res_re),
    .io_res_im(ComplexAdd_io_res_im)
  );
  ComplexSub ComplexSub ( // @[Butterfly.scala 40:22]
    .io_op1_re(ComplexSub_io_op1_re),
    .io_op1_im(ComplexSub_io_op1_im),
    .io_op2_re(ComplexSub_io_op2_re),
    .io_op2_im(ComplexSub_io_op2_im),
    .io_res_re(ComplexSub_io_res_re),
    .io_res_im(ComplexSub_io_res_im)
  );
  assign io_dOut1_re = _T_985_re; // @[FFT.scala 88:12]
  assign io_dOut1_im = _T_985_im; // @[FFT.scala 88:12]
  assign io_dOut2_re = _T_986_re; // @[FFT.scala 89:12]
  assign io_dOut2_im = _T_986_im; // @[FFT.scala 89:12]
  assign io_dout_valid = _T_1498 & _T_2267; // @[FFT.scala 90:17]
  assign Butterfly_io_in1_re = _T_405_re; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in1_im = _T_405_im; // @[Butterfly.scala 90:17]
  assign Butterfly_io_in2_re = io_dIn_re; // @[Butterfly.scala 91:17]
  assign Butterfly_io_in2_im = io_dIn_im; // @[Butterfly.scala 91:17]
  assign Butterfly_io_wn_re = 8'hff == cnt[7:0] ? $signed(-32'shfffb) : $signed(_GEN_255); // @[Butterfly.scala 92:16]
  assign Butterfly_io_wn_im = 8'hff == cnt[7:0] ? $signed(-32'sh324) : $signed(_GEN_1023); // @[Butterfly.scala 92:16]
  assign Switch_io_in1_re = Butterfly_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_io_in1_im = Butterfly_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_io_in2_re = _T_534_re; // @[Butterfly.scala 112:17]
  assign Switch_io_in2_im = _T_534_im; // @[Butterfly.scala 112:17]
  assign Switch_io_sel = cnt[7]; // @[Butterfly.scala 113:17]
  assign Butterfly_1_io_in1_re = _T_670_re; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in1_im = _T_670_im; // @[Butterfly.scala 90:17]
  assign Butterfly_1_io_in2_re = Switch_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_in2_im = Switch_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_1_io_wn_re = 7'h7f == cnt[6:0] ? $signed(-32'shffec) : $signed(_GEN_1919); // @[Butterfly.scala 92:16]
  assign Butterfly_1_io_wn_im = 7'h7f == cnt[6:0] ? $signed(-32'sh648) : $signed(_GEN_2303); // @[Butterfly.scala 92:16]
  assign Switch_1_io_in1_re = Butterfly_1_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in1_im = Butterfly_1_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_1_io_in2_re = _T_735_re; // @[Butterfly.scala 112:17]
  assign Switch_1_io_in2_im = _T_735_im; // @[Butterfly.scala 112:17]
  assign Switch_1_io_sel = cnt[6]; // @[Butterfly.scala 113:17]
  assign Butterfly_2_io_in1_re = _T_807_re; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in1_im = _T_807_im; // @[Butterfly.scala 90:17]
  assign Butterfly_2_io_in2_re = Switch_1_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_in2_im = Switch_1_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_2_io_wn_re = 6'h3f == cnt[5:0] ? $signed(-32'shffb1) : $signed(_GEN_2751); // @[Butterfly.scala 92:16]
  assign Butterfly_2_io_wn_im = 6'h3f == cnt[5:0] ? $signed(-32'shc90) : $signed(_GEN_2943); // @[Butterfly.scala 92:16]
  assign Switch_2_io_in1_re = Butterfly_2_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in1_im = Butterfly_2_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_2_io_in2_re = _T_840_re; // @[Butterfly.scala 112:17]
  assign Switch_2_io_in2_im = _T_840_im; // @[Butterfly.scala 112:17]
  assign Switch_2_io_sel = cnt[5]; // @[Butterfly.scala 113:17]
  assign Butterfly_3_io_in1_re = _T_880_re; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in1_im = _T_880_im; // @[Butterfly.scala 90:17]
  assign Butterfly_3_io_in2_re = Switch_2_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_in2_im = Switch_2_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_3_io_wn_re = 5'h1f == cnt[4:0] ? $signed(-32'shfec4) : $signed(_GEN_3167); // @[Butterfly.scala 92:16]
  assign Butterfly_3_io_wn_im = 5'h1f == cnt[4:0] ? $signed(-32'sh1918) : $signed(_GEN_3263); // @[Butterfly.scala 92:16]
  assign Switch_3_io_in1_re = Butterfly_3_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in1_im = Butterfly_3_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_3_io_in2_re = _T_897_re; // @[Butterfly.scala 112:17]
  assign Switch_3_io_in2_im = _T_897_im; // @[Butterfly.scala 112:17]
  assign Switch_3_io_sel = cnt[4]; // @[Butterfly.scala 113:17]
  assign Butterfly_4_io_in1_re = _T_921_re; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in1_im = _T_921_im; // @[Butterfly.scala 90:17]
  assign Butterfly_4_io_in2_re = Switch_3_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_in2_im = Switch_3_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_4_io_wn_re = 4'hf == cnt[3:0] ? $signed(-32'shfb15) : $signed(_GEN_3375); // @[Butterfly.scala 92:16]
  assign Butterfly_4_io_wn_im = 4'hf == cnt[3:0] ? $signed(-32'sh31f1) : $signed(_GEN_3423); // @[Butterfly.scala 92:16]
  assign Switch_4_io_in1_re = Butterfly_4_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in1_im = Butterfly_4_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_4_io_in2_re = _T_930_re; // @[Butterfly.scala 112:17]
  assign Switch_4_io_in2_im = _T_930_im; // @[Butterfly.scala 112:17]
  assign Switch_4_io_sel = cnt[3]; // @[Butterfly.scala 113:17]
  assign Butterfly_5_io_in1_re = _T_946_re; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in1_im = _T_946_im; // @[Butterfly.scala 90:17]
  assign Butterfly_5_io_in2_re = Switch_4_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_in2_im = Switch_4_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_5_io_wn_re = 3'h7 == cnt[2:0] ? $signed(-32'shec83) : $signed(_GEN_3479); // @[Butterfly.scala 92:16]
  assign Butterfly_5_io_wn_im = 3'h7 == cnt[2:0] ? $signed(-32'sh61f8) : $signed(_GEN_3503); // @[Butterfly.scala 92:16]
  assign Switch_5_io_in1_re = Butterfly_5_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in1_im = Butterfly_5_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_5_io_in2_re = _T_951_re; // @[Butterfly.scala 112:17]
  assign Switch_5_io_in2_im = _T_951_im; // @[Butterfly.scala 112:17]
  assign Switch_5_io_sel = cnt[2]; // @[Butterfly.scala 113:17]
  assign Butterfly_6_io_in1_re = _T_963_re; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in1_im = _T_963_im; // @[Butterfly.scala 90:17]
  assign Butterfly_6_io_in2_re = Switch_5_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_in2_im = Switch_5_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_6_io_wn_re = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_3531); // @[Butterfly.scala 92:16]
  assign Butterfly_6_io_wn_im = 2'h3 == cnt[1:0] ? $signed(-32'shb505) : $signed(_GEN_3543); // @[Butterfly.scala 92:16]
  assign Switch_6_io_in1_re = Butterfly_6_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in1_im = Butterfly_6_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_6_io_in2_re = _T_966_re; // @[Butterfly.scala 112:17]
  assign Switch_6_io_in2_im = _T_966_im; // @[Butterfly.scala 112:17]
  assign Switch_6_io_sel = cnt[1]; // @[Butterfly.scala 113:17]
  assign Butterfly_7_io_in1_re = _T_976_re; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in1_im = _T_976_im; // @[Butterfly.scala 90:17]
  assign Butterfly_7_io_in2_re = Switch_6_io_out2_re; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_in2_im = Switch_6_io_out2_im; // @[Butterfly.scala 91:17]
  assign Butterfly_7_io_wn_re = cnt[0] ? $signed(32'sh0) : $signed(32'sh10000); // @[Butterfly.scala 92:16]
  assign Butterfly_7_io_wn_im = cnt[0] ? $signed(-32'sh10000) : $signed(32'sh0); // @[Butterfly.scala 92:16]
  assign Switch_7_io_in1_re = Butterfly_7_io_out1_re; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in1_im = Butterfly_7_io_out1_im; // @[Butterfly.scala 111:17]
  assign Switch_7_io_in2_re = _T_978_re; // @[Butterfly.scala 112:17]
  assign Switch_7_io_in2_im = _T_978_im; // @[Butterfly.scala 112:17]
  assign Switch_7_io_sel = cnt[0]; // @[Butterfly.scala 113:17]
  assign ComplexAdd_io_op1_re = out1D1_re; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op1_im = out1D1_im; // @[Butterfly.scala 27:17]
  assign ComplexAdd_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 28:17]
  assign ComplexAdd_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 28:17]
  assign ComplexSub_io_op1_re = out1D1_re; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op1_im = out1D1_im; // @[Butterfly.scala 41:17]
  assign ComplexSub_io_op2_re = Switch_7_io_out2_re; // @[Butterfly.scala 42:17]
  assign ComplexSub_io_op2_im = Switch_7_io_out2_im; // @[Butterfly.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  _T_150_re = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_150_im = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  _T_151_re = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  _T_151_im = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  _T_152_re = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  _T_152_im = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _T_153_re = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _T_153_im = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  _T_154_re = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  _T_154_im = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  _T_155_re = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _T_155_im = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  _T_156_re = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  _T_156_im = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  _T_157_re = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  _T_157_im = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  _T_158_re = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  _T_158_im = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  _T_159_re = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  _T_159_im = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  _T_160_re = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  _T_160_im = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  _T_161_re = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  _T_161_im = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  _T_162_re = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  _T_162_im = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  _T_163_re = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  _T_163_im = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  _T_164_re = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  _T_164_im = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  _T_165_re = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  _T_165_im = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  _T_166_re = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  _T_166_im = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  _T_167_re = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  _T_167_im = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  _T_168_re = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  _T_168_im = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  _T_169_re = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  _T_169_im = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  _T_170_re = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  _T_170_im = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  _T_171_re = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  _T_171_im = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  _T_172_re = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  _T_172_im = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  _T_173_re = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  _T_173_im = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  _T_174_re = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  _T_174_im = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  _T_175_re = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  _T_175_im = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  _T_176_re = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  _T_176_im = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  _T_177_re = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  _T_177_im = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  _T_178_re = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  _T_178_im = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  _T_179_re = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  _T_179_im = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  _T_180_re = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  _T_180_im = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  _T_181_re = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  _T_181_im = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  _T_182_re = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  _T_182_im = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  _T_183_re = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  _T_183_im = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  _T_184_re = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  _T_184_im = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  _T_185_re = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  _T_185_im = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  _T_186_re = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  _T_186_im = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  _T_187_re = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  _T_187_im = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  _T_188_re = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  _T_188_im = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  _T_189_re = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  _T_189_im = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  _T_190_re = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  _T_190_im = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  _T_191_re = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  _T_191_im = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  _T_192_re = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  _T_192_im = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  _T_193_re = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  _T_193_im = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  _T_194_re = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  _T_194_im = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  _T_195_re = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  _T_195_im = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  _T_196_re = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  _T_196_im = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  _T_197_re = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  _T_197_im = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  _T_198_re = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  _T_198_im = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  _T_199_re = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  _T_199_im = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  _T_200_re = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  _T_200_im = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  _T_201_re = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  _T_201_im = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  _T_202_re = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  _T_202_im = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  _T_203_re = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  _T_203_im = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  _T_204_re = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  _T_204_im = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  _T_205_re = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  _T_205_im = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  _T_206_re = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  _T_206_im = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  _T_207_re = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  _T_207_im = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  _T_208_re = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  _T_208_im = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  _T_209_re = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  _T_209_im = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  _T_210_re = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  _T_210_im = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  _T_211_re = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  _T_211_im = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  _T_212_re = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  _T_212_im = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  _T_213_re = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  _T_213_im = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  _T_214_re = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  _T_214_im = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  _T_215_re = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  _T_215_im = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  _T_216_re = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  _T_216_im = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  _T_217_re = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  _T_217_im = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  _T_218_re = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  _T_218_im = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  _T_219_re = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  _T_219_im = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  _T_220_re = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  _T_220_im = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  _T_221_re = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  _T_221_im = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  _T_222_re = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  _T_222_im = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  _T_223_re = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  _T_223_im = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  _T_224_re = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  _T_224_im = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  _T_225_re = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  _T_225_im = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  _T_226_re = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  _T_226_im = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  _T_227_re = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  _T_227_im = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  _T_228_re = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  _T_228_im = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  _T_229_re = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  _T_229_im = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  _T_230_re = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  _T_230_im = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  _T_231_re = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  _T_231_im = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  _T_232_re = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  _T_232_im = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  _T_233_re = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  _T_233_im = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  _T_234_re = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  _T_234_im = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  _T_235_re = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  _T_235_im = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  _T_236_re = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  _T_236_im = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  _T_237_re = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  _T_237_im = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  _T_238_re = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  _T_238_im = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  _T_239_re = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  _T_239_im = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  _T_240_re = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  _T_240_im = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  _T_241_re = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  _T_241_im = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  _T_242_re = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  _T_242_im = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  _T_243_re = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  _T_243_im = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  _T_244_re = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  _T_244_im = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  _T_245_re = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  _T_245_im = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  _T_246_re = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  _T_246_im = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  _T_247_re = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  _T_247_im = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  _T_248_re = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  _T_248_im = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  _T_249_re = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  _T_249_im = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  _T_250_re = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  _T_250_im = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  _T_251_re = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  _T_251_im = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  _T_252_re = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  _T_252_im = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  _T_253_re = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  _T_253_im = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  _T_254_re = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  _T_254_im = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  _T_255_re = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  _T_255_im = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  _T_256_re = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  _T_256_im = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  _T_257_re = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  _T_257_im = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  _T_258_re = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  _T_258_im = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  _T_259_re = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  _T_259_im = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  _T_260_re = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  _T_260_im = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  _T_261_re = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  _T_261_im = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  _T_262_re = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  _T_262_im = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  _T_263_re = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  _T_263_im = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  _T_264_re = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  _T_264_im = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  _T_265_re = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  _T_265_im = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  _T_266_re = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  _T_266_im = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  _T_267_re = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  _T_267_im = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  _T_268_re = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  _T_268_im = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  _T_269_re = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  _T_269_im = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  _T_270_re = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  _T_270_im = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  _T_271_re = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  _T_271_im = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  _T_272_re = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  _T_272_im = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  _T_273_re = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  _T_273_im = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  _T_274_re = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  _T_274_im = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  _T_275_re = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  _T_275_im = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  _T_276_re = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  _T_276_im = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  _T_277_re = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  _T_277_im = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  _T_278_re = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  _T_278_im = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  _T_279_re = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  _T_279_im = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  _T_280_re = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  _T_280_im = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  _T_281_re = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  _T_281_im = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  _T_282_re = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  _T_282_im = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  _T_283_re = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  _T_283_im = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  _T_284_re = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  _T_284_im = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  _T_285_re = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  _T_285_im = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  _T_286_re = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  _T_286_im = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  _T_287_re = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  _T_287_im = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  _T_288_re = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  _T_288_im = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  _T_289_re = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  _T_289_im = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  _T_290_re = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  _T_290_im = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  _T_291_re = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  _T_291_im = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  _T_292_re = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  _T_292_im = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  _T_293_re = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  _T_293_im = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  _T_294_re = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  _T_294_im = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  _T_295_re = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  _T_295_im = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  _T_296_re = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  _T_296_im = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  _T_297_re = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  _T_297_im = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  _T_298_re = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  _T_298_im = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  _T_299_re = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  _T_299_im = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  _T_300_re = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  _T_300_im = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  _T_301_re = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  _T_301_im = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  _T_302_re = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  _T_302_im = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  _T_303_re = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  _T_303_im = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  _T_304_re = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  _T_304_im = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  _T_305_re = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  _T_305_im = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  _T_306_re = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  _T_306_im = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  _T_307_re = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  _T_307_im = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  _T_308_re = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  _T_308_im = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  _T_309_re = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  _T_309_im = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  _T_310_re = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  _T_310_im = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  _T_311_re = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  _T_311_im = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  _T_312_re = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  _T_312_im = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  _T_313_re = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  _T_313_im = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  _T_314_re = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  _T_314_im = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  _T_315_re = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  _T_315_im = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  _T_316_re = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  _T_316_im = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  _T_317_re = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  _T_317_im = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  _T_318_re = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  _T_318_im = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  _T_319_re = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  _T_319_im = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  _T_320_re = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  _T_320_im = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  _T_321_re = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  _T_321_im = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  _T_322_re = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  _T_322_im = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  _T_323_re = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  _T_323_im = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  _T_324_re = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  _T_324_im = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  _T_325_re = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  _T_325_im = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  _T_326_re = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  _T_326_im = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  _T_327_re = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  _T_327_im = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  _T_328_re = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  _T_328_im = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  _T_329_re = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  _T_329_im = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  _T_330_re = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  _T_330_im = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  _T_331_re = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  _T_331_im = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  _T_332_re = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  _T_332_im = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  _T_333_re = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  _T_333_im = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  _T_334_re = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  _T_334_im = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  _T_335_re = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  _T_335_im = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  _T_336_re = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  _T_336_im = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  _T_337_re = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  _T_337_im = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  _T_338_re = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  _T_338_im = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  _T_339_re = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  _T_339_im = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  _T_340_re = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  _T_340_im = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  _T_341_re = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  _T_341_im = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  _T_342_re = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  _T_342_im = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  _T_343_re = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  _T_343_im = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  _T_344_re = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  _T_344_im = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  _T_345_re = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  _T_345_im = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  _T_346_re = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  _T_346_im = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  _T_347_re = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  _T_347_im = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  _T_348_re = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  _T_348_im = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  _T_349_re = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  _T_349_im = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  _T_350_re = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  _T_350_im = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  _T_351_re = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  _T_351_im = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  _T_352_re = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  _T_352_im = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  _T_353_re = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  _T_353_im = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  _T_354_re = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  _T_354_im = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  _T_355_re = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  _T_355_im = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  _T_356_re = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  _T_356_im = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  _T_357_re = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  _T_357_im = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  _T_358_re = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  _T_358_im = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  _T_359_re = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  _T_359_im = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  _T_360_re = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  _T_360_im = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  _T_361_re = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  _T_361_im = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  _T_362_re = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  _T_362_im = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  _T_363_re = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  _T_363_im = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  _T_364_re = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  _T_364_im = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  _T_365_re = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  _T_365_im = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  _T_366_re = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  _T_366_im = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  _T_367_re = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  _T_367_im = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  _T_368_re = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  _T_368_im = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  _T_369_re = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  _T_369_im = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  _T_370_re = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  _T_370_im = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  _T_371_re = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  _T_371_im = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  _T_372_re = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  _T_372_im = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  _T_373_re = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  _T_373_im = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  _T_374_re = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  _T_374_im = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  _T_375_re = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  _T_375_im = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  _T_376_re = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  _T_376_im = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  _T_377_re = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  _T_377_im = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  _T_378_re = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  _T_378_im = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  _T_379_re = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  _T_379_im = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  _T_380_re = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  _T_380_im = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  _T_381_re = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  _T_381_im = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  _T_382_re = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  _T_382_im = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  _T_383_re = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  _T_383_im = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  _T_384_re = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  _T_384_im = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  _T_385_re = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  _T_385_im = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  _T_386_re = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  _T_386_im = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  _T_387_re = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  _T_387_im = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  _T_388_re = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  _T_388_im = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  _T_389_re = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  _T_389_im = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  _T_390_re = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  _T_390_im = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  _T_391_re = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  _T_391_im = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  _T_392_re = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  _T_392_im = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  _T_393_re = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  _T_393_im = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  _T_394_re = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  _T_394_im = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  _T_395_re = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  _T_395_im = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  _T_396_re = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  _T_396_im = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  _T_397_re = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  _T_397_im = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  _T_398_re = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  _T_398_im = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  _T_399_re = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  _T_399_im = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  _T_400_re = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  _T_400_im = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  _T_401_re = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  _T_401_im = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  _T_402_re = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  _T_402_im = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  _T_403_re = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  _T_403_im = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  _T_404_re = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  _T_404_im = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  _T_405_re = _RAND_511[31:0];
  _RAND_512 = {1{`RANDOM}};
  _T_405_im = _RAND_512[31:0];
  _RAND_513 = {1{`RANDOM}};
  _T_407_re = _RAND_513[31:0];
  _RAND_514 = {1{`RANDOM}};
  _T_407_im = _RAND_514[31:0];
  _RAND_515 = {1{`RANDOM}};
  _T_408_re = _RAND_515[31:0];
  _RAND_516 = {1{`RANDOM}};
  _T_408_im = _RAND_516[31:0];
  _RAND_517 = {1{`RANDOM}};
  _T_409_re = _RAND_517[31:0];
  _RAND_518 = {1{`RANDOM}};
  _T_409_im = _RAND_518[31:0];
  _RAND_519 = {1{`RANDOM}};
  _T_410_re = _RAND_519[31:0];
  _RAND_520 = {1{`RANDOM}};
  _T_410_im = _RAND_520[31:0];
  _RAND_521 = {1{`RANDOM}};
  _T_411_re = _RAND_521[31:0];
  _RAND_522 = {1{`RANDOM}};
  _T_411_im = _RAND_522[31:0];
  _RAND_523 = {1{`RANDOM}};
  _T_412_re = _RAND_523[31:0];
  _RAND_524 = {1{`RANDOM}};
  _T_412_im = _RAND_524[31:0];
  _RAND_525 = {1{`RANDOM}};
  _T_413_re = _RAND_525[31:0];
  _RAND_526 = {1{`RANDOM}};
  _T_413_im = _RAND_526[31:0];
  _RAND_527 = {1{`RANDOM}};
  _T_414_re = _RAND_527[31:0];
  _RAND_528 = {1{`RANDOM}};
  _T_414_im = _RAND_528[31:0];
  _RAND_529 = {1{`RANDOM}};
  _T_415_re = _RAND_529[31:0];
  _RAND_530 = {1{`RANDOM}};
  _T_415_im = _RAND_530[31:0];
  _RAND_531 = {1{`RANDOM}};
  _T_416_re = _RAND_531[31:0];
  _RAND_532 = {1{`RANDOM}};
  _T_416_im = _RAND_532[31:0];
  _RAND_533 = {1{`RANDOM}};
  _T_417_re = _RAND_533[31:0];
  _RAND_534 = {1{`RANDOM}};
  _T_417_im = _RAND_534[31:0];
  _RAND_535 = {1{`RANDOM}};
  _T_418_re = _RAND_535[31:0];
  _RAND_536 = {1{`RANDOM}};
  _T_418_im = _RAND_536[31:0];
  _RAND_537 = {1{`RANDOM}};
  _T_419_re = _RAND_537[31:0];
  _RAND_538 = {1{`RANDOM}};
  _T_419_im = _RAND_538[31:0];
  _RAND_539 = {1{`RANDOM}};
  _T_420_re = _RAND_539[31:0];
  _RAND_540 = {1{`RANDOM}};
  _T_420_im = _RAND_540[31:0];
  _RAND_541 = {1{`RANDOM}};
  _T_421_re = _RAND_541[31:0];
  _RAND_542 = {1{`RANDOM}};
  _T_421_im = _RAND_542[31:0];
  _RAND_543 = {1{`RANDOM}};
  _T_422_re = _RAND_543[31:0];
  _RAND_544 = {1{`RANDOM}};
  _T_422_im = _RAND_544[31:0];
  _RAND_545 = {1{`RANDOM}};
  _T_423_re = _RAND_545[31:0];
  _RAND_546 = {1{`RANDOM}};
  _T_423_im = _RAND_546[31:0];
  _RAND_547 = {1{`RANDOM}};
  _T_424_re = _RAND_547[31:0];
  _RAND_548 = {1{`RANDOM}};
  _T_424_im = _RAND_548[31:0];
  _RAND_549 = {1{`RANDOM}};
  _T_425_re = _RAND_549[31:0];
  _RAND_550 = {1{`RANDOM}};
  _T_425_im = _RAND_550[31:0];
  _RAND_551 = {1{`RANDOM}};
  _T_426_re = _RAND_551[31:0];
  _RAND_552 = {1{`RANDOM}};
  _T_426_im = _RAND_552[31:0];
  _RAND_553 = {1{`RANDOM}};
  _T_427_re = _RAND_553[31:0];
  _RAND_554 = {1{`RANDOM}};
  _T_427_im = _RAND_554[31:0];
  _RAND_555 = {1{`RANDOM}};
  _T_428_re = _RAND_555[31:0];
  _RAND_556 = {1{`RANDOM}};
  _T_428_im = _RAND_556[31:0];
  _RAND_557 = {1{`RANDOM}};
  _T_429_re = _RAND_557[31:0];
  _RAND_558 = {1{`RANDOM}};
  _T_429_im = _RAND_558[31:0];
  _RAND_559 = {1{`RANDOM}};
  _T_430_re = _RAND_559[31:0];
  _RAND_560 = {1{`RANDOM}};
  _T_430_im = _RAND_560[31:0];
  _RAND_561 = {1{`RANDOM}};
  _T_431_re = _RAND_561[31:0];
  _RAND_562 = {1{`RANDOM}};
  _T_431_im = _RAND_562[31:0];
  _RAND_563 = {1{`RANDOM}};
  _T_432_re = _RAND_563[31:0];
  _RAND_564 = {1{`RANDOM}};
  _T_432_im = _RAND_564[31:0];
  _RAND_565 = {1{`RANDOM}};
  _T_433_re = _RAND_565[31:0];
  _RAND_566 = {1{`RANDOM}};
  _T_433_im = _RAND_566[31:0];
  _RAND_567 = {1{`RANDOM}};
  _T_434_re = _RAND_567[31:0];
  _RAND_568 = {1{`RANDOM}};
  _T_434_im = _RAND_568[31:0];
  _RAND_569 = {1{`RANDOM}};
  _T_435_re = _RAND_569[31:0];
  _RAND_570 = {1{`RANDOM}};
  _T_435_im = _RAND_570[31:0];
  _RAND_571 = {1{`RANDOM}};
  _T_436_re = _RAND_571[31:0];
  _RAND_572 = {1{`RANDOM}};
  _T_436_im = _RAND_572[31:0];
  _RAND_573 = {1{`RANDOM}};
  _T_437_re = _RAND_573[31:0];
  _RAND_574 = {1{`RANDOM}};
  _T_437_im = _RAND_574[31:0];
  _RAND_575 = {1{`RANDOM}};
  _T_438_re = _RAND_575[31:0];
  _RAND_576 = {1{`RANDOM}};
  _T_438_im = _RAND_576[31:0];
  _RAND_577 = {1{`RANDOM}};
  _T_439_re = _RAND_577[31:0];
  _RAND_578 = {1{`RANDOM}};
  _T_439_im = _RAND_578[31:0];
  _RAND_579 = {1{`RANDOM}};
  _T_440_re = _RAND_579[31:0];
  _RAND_580 = {1{`RANDOM}};
  _T_440_im = _RAND_580[31:0];
  _RAND_581 = {1{`RANDOM}};
  _T_441_re = _RAND_581[31:0];
  _RAND_582 = {1{`RANDOM}};
  _T_441_im = _RAND_582[31:0];
  _RAND_583 = {1{`RANDOM}};
  _T_442_re = _RAND_583[31:0];
  _RAND_584 = {1{`RANDOM}};
  _T_442_im = _RAND_584[31:0];
  _RAND_585 = {1{`RANDOM}};
  _T_443_re = _RAND_585[31:0];
  _RAND_586 = {1{`RANDOM}};
  _T_443_im = _RAND_586[31:0];
  _RAND_587 = {1{`RANDOM}};
  _T_444_re = _RAND_587[31:0];
  _RAND_588 = {1{`RANDOM}};
  _T_444_im = _RAND_588[31:0];
  _RAND_589 = {1{`RANDOM}};
  _T_445_re = _RAND_589[31:0];
  _RAND_590 = {1{`RANDOM}};
  _T_445_im = _RAND_590[31:0];
  _RAND_591 = {1{`RANDOM}};
  _T_446_re = _RAND_591[31:0];
  _RAND_592 = {1{`RANDOM}};
  _T_446_im = _RAND_592[31:0];
  _RAND_593 = {1{`RANDOM}};
  _T_447_re = _RAND_593[31:0];
  _RAND_594 = {1{`RANDOM}};
  _T_447_im = _RAND_594[31:0];
  _RAND_595 = {1{`RANDOM}};
  _T_448_re = _RAND_595[31:0];
  _RAND_596 = {1{`RANDOM}};
  _T_448_im = _RAND_596[31:0];
  _RAND_597 = {1{`RANDOM}};
  _T_449_re = _RAND_597[31:0];
  _RAND_598 = {1{`RANDOM}};
  _T_449_im = _RAND_598[31:0];
  _RAND_599 = {1{`RANDOM}};
  _T_450_re = _RAND_599[31:0];
  _RAND_600 = {1{`RANDOM}};
  _T_450_im = _RAND_600[31:0];
  _RAND_601 = {1{`RANDOM}};
  _T_451_re = _RAND_601[31:0];
  _RAND_602 = {1{`RANDOM}};
  _T_451_im = _RAND_602[31:0];
  _RAND_603 = {1{`RANDOM}};
  _T_452_re = _RAND_603[31:0];
  _RAND_604 = {1{`RANDOM}};
  _T_452_im = _RAND_604[31:0];
  _RAND_605 = {1{`RANDOM}};
  _T_453_re = _RAND_605[31:0];
  _RAND_606 = {1{`RANDOM}};
  _T_453_im = _RAND_606[31:0];
  _RAND_607 = {1{`RANDOM}};
  _T_454_re = _RAND_607[31:0];
  _RAND_608 = {1{`RANDOM}};
  _T_454_im = _RAND_608[31:0];
  _RAND_609 = {1{`RANDOM}};
  _T_455_re = _RAND_609[31:0];
  _RAND_610 = {1{`RANDOM}};
  _T_455_im = _RAND_610[31:0];
  _RAND_611 = {1{`RANDOM}};
  _T_456_re = _RAND_611[31:0];
  _RAND_612 = {1{`RANDOM}};
  _T_456_im = _RAND_612[31:0];
  _RAND_613 = {1{`RANDOM}};
  _T_457_re = _RAND_613[31:0];
  _RAND_614 = {1{`RANDOM}};
  _T_457_im = _RAND_614[31:0];
  _RAND_615 = {1{`RANDOM}};
  _T_458_re = _RAND_615[31:0];
  _RAND_616 = {1{`RANDOM}};
  _T_458_im = _RAND_616[31:0];
  _RAND_617 = {1{`RANDOM}};
  _T_459_re = _RAND_617[31:0];
  _RAND_618 = {1{`RANDOM}};
  _T_459_im = _RAND_618[31:0];
  _RAND_619 = {1{`RANDOM}};
  _T_460_re = _RAND_619[31:0];
  _RAND_620 = {1{`RANDOM}};
  _T_460_im = _RAND_620[31:0];
  _RAND_621 = {1{`RANDOM}};
  _T_461_re = _RAND_621[31:0];
  _RAND_622 = {1{`RANDOM}};
  _T_461_im = _RAND_622[31:0];
  _RAND_623 = {1{`RANDOM}};
  _T_462_re = _RAND_623[31:0];
  _RAND_624 = {1{`RANDOM}};
  _T_462_im = _RAND_624[31:0];
  _RAND_625 = {1{`RANDOM}};
  _T_463_re = _RAND_625[31:0];
  _RAND_626 = {1{`RANDOM}};
  _T_463_im = _RAND_626[31:0];
  _RAND_627 = {1{`RANDOM}};
  _T_464_re = _RAND_627[31:0];
  _RAND_628 = {1{`RANDOM}};
  _T_464_im = _RAND_628[31:0];
  _RAND_629 = {1{`RANDOM}};
  _T_465_re = _RAND_629[31:0];
  _RAND_630 = {1{`RANDOM}};
  _T_465_im = _RAND_630[31:0];
  _RAND_631 = {1{`RANDOM}};
  _T_466_re = _RAND_631[31:0];
  _RAND_632 = {1{`RANDOM}};
  _T_466_im = _RAND_632[31:0];
  _RAND_633 = {1{`RANDOM}};
  _T_467_re = _RAND_633[31:0];
  _RAND_634 = {1{`RANDOM}};
  _T_467_im = _RAND_634[31:0];
  _RAND_635 = {1{`RANDOM}};
  _T_468_re = _RAND_635[31:0];
  _RAND_636 = {1{`RANDOM}};
  _T_468_im = _RAND_636[31:0];
  _RAND_637 = {1{`RANDOM}};
  _T_469_re = _RAND_637[31:0];
  _RAND_638 = {1{`RANDOM}};
  _T_469_im = _RAND_638[31:0];
  _RAND_639 = {1{`RANDOM}};
  _T_470_re = _RAND_639[31:0];
  _RAND_640 = {1{`RANDOM}};
  _T_470_im = _RAND_640[31:0];
  _RAND_641 = {1{`RANDOM}};
  _T_471_re = _RAND_641[31:0];
  _RAND_642 = {1{`RANDOM}};
  _T_471_im = _RAND_642[31:0];
  _RAND_643 = {1{`RANDOM}};
  _T_472_re = _RAND_643[31:0];
  _RAND_644 = {1{`RANDOM}};
  _T_472_im = _RAND_644[31:0];
  _RAND_645 = {1{`RANDOM}};
  _T_473_re = _RAND_645[31:0];
  _RAND_646 = {1{`RANDOM}};
  _T_473_im = _RAND_646[31:0];
  _RAND_647 = {1{`RANDOM}};
  _T_474_re = _RAND_647[31:0];
  _RAND_648 = {1{`RANDOM}};
  _T_474_im = _RAND_648[31:0];
  _RAND_649 = {1{`RANDOM}};
  _T_475_re = _RAND_649[31:0];
  _RAND_650 = {1{`RANDOM}};
  _T_475_im = _RAND_650[31:0];
  _RAND_651 = {1{`RANDOM}};
  _T_476_re = _RAND_651[31:0];
  _RAND_652 = {1{`RANDOM}};
  _T_476_im = _RAND_652[31:0];
  _RAND_653 = {1{`RANDOM}};
  _T_477_re = _RAND_653[31:0];
  _RAND_654 = {1{`RANDOM}};
  _T_477_im = _RAND_654[31:0];
  _RAND_655 = {1{`RANDOM}};
  _T_478_re = _RAND_655[31:0];
  _RAND_656 = {1{`RANDOM}};
  _T_478_im = _RAND_656[31:0];
  _RAND_657 = {1{`RANDOM}};
  _T_479_re = _RAND_657[31:0];
  _RAND_658 = {1{`RANDOM}};
  _T_479_im = _RAND_658[31:0];
  _RAND_659 = {1{`RANDOM}};
  _T_480_re = _RAND_659[31:0];
  _RAND_660 = {1{`RANDOM}};
  _T_480_im = _RAND_660[31:0];
  _RAND_661 = {1{`RANDOM}};
  _T_481_re = _RAND_661[31:0];
  _RAND_662 = {1{`RANDOM}};
  _T_481_im = _RAND_662[31:0];
  _RAND_663 = {1{`RANDOM}};
  _T_482_re = _RAND_663[31:0];
  _RAND_664 = {1{`RANDOM}};
  _T_482_im = _RAND_664[31:0];
  _RAND_665 = {1{`RANDOM}};
  _T_483_re = _RAND_665[31:0];
  _RAND_666 = {1{`RANDOM}};
  _T_483_im = _RAND_666[31:0];
  _RAND_667 = {1{`RANDOM}};
  _T_484_re = _RAND_667[31:0];
  _RAND_668 = {1{`RANDOM}};
  _T_484_im = _RAND_668[31:0];
  _RAND_669 = {1{`RANDOM}};
  _T_485_re = _RAND_669[31:0];
  _RAND_670 = {1{`RANDOM}};
  _T_485_im = _RAND_670[31:0];
  _RAND_671 = {1{`RANDOM}};
  _T_486_re = _RAND_671[31:0];
  _RAND_672 = {1{`RANDOM}};
  _T_486_im = _RAND_672[31:0];
  _RAND_673 = {1{`RANDOM}};
  _T_487_re = _RAND_673[31:0];
  _RAND_674 = {1{`RANDOM}};
  _T_487_im = _RAND_674[31:0];
  _RAND_675 = {1{`RANDOM}};
  _T_488_re = _RAND_675[31:0];
  _RAND_676 = {1{`RANDOM}};
  _T_488_im = _RAND_676[31:0];
  _RAND_677 = {1{`RANDOM}};
  _T_489_re = _RAND_677[31:0];
  _RAND_678 = {1{`RANDOM}};
  _T_489_im = _RAND_678[31:0];
  _RAND_679 = {1{`RANDOM}};
  _T_490_re = _RAND_679[31:0];
  _RAND_680 = {1{`RANDOM}};
  _T_490_im = _RAND_680[31:0];
  _RAND_681 = {1{`RANDOM}};
  _T_491_re = _RAND_681[31:0];
  _RAND_682 = {1{`RANDOM}};
  _T_491_im = _RAND_682[31:0];
  _RAND_683 = {1{`RANDOM}};
  _T_492_re = _RAND_683[31:0];
  _RAND_684 = {1{`RANDOM}};
  _T_492_im = _RAND_684[31:0];
  _RAND_685 = {1{`RANDOM}};
  _T_493_re = _RAND_685[31:0];
  _RAND_686 = {1{`RANDOM}};
  _T_493_im = _RAND_686[31:0];
  _RAND_687 = {1{`RANDOM}};
  _T_494_re = _RAND_687[31:0];
  _RAND_688 = {1{`RANDOM}};
  _T_494_im = _RAND_688[31:0];
  _RAND_689 = {1{`RANDOM}};
  _T_495_re = _RAND_689[31:0];
  _RAND_690 = {1{`RANDOM}};
  _T_495_im = _RAND_690[31:0];
  _RAND_691 = {1{`RANDOM}};
  _T_496_re = _RAND_691[31:0];
  _RAND_692 = {1{`RANDOM}};
  _T_496_im = _RAND_692[31:0];
  _RAND_693 = {1{`RANDOM}};
  _T_497_re = _RAND_693[31:0];
  _RAND_694 = {1{`RANDOM}};
  _T_497_im = _RAND_694[31:0];
  _RAND_695 = {1{`RANDOM}};
  _T_498_re = _RAND_695[31:0];
  _RAND_696 = {1{`RANDOM}};
  _T_498_im = _RAND_696[31:0];
  _RAND_697 = {1{`RANDOM}};
  _T_499_re = _RAND_697[31:0];
  _RAND_698 = {1{`RANDOM}};
  _T_499_im = _RAND_698[31:0];
  _RAND_699 = {1{`RANDOM}};
  _T_500_re = _RAND_699[31:0];
  _RAND_700 = {1{`RANDOM}};
  _T_500_im = _RAND_700[31:0];
  _RAND_701 = {1{`RANDOM}};
  _T_501_re = _RAND_701[31:0];
  _RAND_702 = {1{`RANDOM}};
  _T_501_im = _RAND_702[31:0];
  _RAND_703 = {1{`RANDOM}};
  _T_502_re = _RAND_703[31:0];
  _RAND_704 = {1{`RANDOM}};
  _T_502_im = _RAND_704[31:0];
  _RAND_705 = {1{`RANDOM}};
  _T_503_re = _RAND_705[31:0];
  _RAND_706 = {1{`RANDOM}};
  _T_503_im = _RAND_706[31:0];
  _RAND_707 = {1{`RANDOM}};
  _T_504_re = _RAND_707[31:0];
  _RAND_708 = {1{`RANDOM}};
  _T_504_im = _RAND_708[31:0];
  _RAND_709 = {1{`RANDOM}};
  _T_505_re = _RAND_709[31:0];
  _RAND_710 = {1{`RANDOM}};
  _T_505_im = _RAND_710[31:0];
  _RAND_711 = {1{`RANDOM}};
  _T_506_re = _RAND_711[31:0];
  _RAND_712 = {1{`RANDOM}};
  _T_506_im = _RAND_712[31:0];
  _RAND_713 = {1{`RANDOM}};
  _T_507_re = _RAND_713[31:0];
  _RAND_714 = {1{`RANDOM}};
  _T_507_im = _RAND_714[31:0];
  _RAND_715 = {1{`RANDOM}};
  _T_508_re = _RAND_715[31:0];
  _RAND_716 = {1{`RANDOM}};
  _T_508_im = _RAND_716[31:0];
  _RAND_717 = {1{`RANDOM}};
  _T_509_re = _RAND_717[31:0];
  _RAND_718 = {1{`RANDOM}};
  _T_509_im = _RAND_718[31:0];
  _RAND_719 = {1{`RANDOM}};
  _T_510_re = _RAND_719[31:0];
  _RAND_720 = {1{`RANDOM}};
  _T_510_im = _RAND_720[31:0];
  _RAND_721 = {1{`RANDOM}};
  _T_511_re = _RAND_721[31:0];
  _RAND_722 = {1{`RANDOM}};
  _T_511_im = _RAND_722[31:0];
  _RAND_723 = {1{`RANDOM}};
  _T_512_re = _RAND_723[31:0];
  _RAND_724 = {1{`RANDOM}};
  _T_512_im = _RAND_724[31:0];
  _RAND_725 = {1{`RANDOM}};
  _T_513_re = _RAND_725[31:0];
  _RAND_726 = {1{`RANDOM}};
  _T_513_im = _RAND_726[31:0];
  _RAND_727 = {1{`RANDOM}};
  _T_514_re = _RAND_727[31:0];
  _RAND_728 = {1{`RANDOM}};
  _T_514_im = _RAND_728[31:0];
  _RAND_729 = {1{`RANDOM}};
  _T_515_re = _RAND_729[31:0];
  _RAND_730 = {1{`RANDOM}};
  _T_515_im = _RAND_730[31:0];
  _RAND_731 = {1{`RANDOM}};
  _T_516_re = _RAND_731[31:0];
  _RAND_732 = {1{`RANDOM}};
  _T_516_im = _RAND_732[31:0];
  _RAND_733 = {1{`RANDOM}};
  _T_517_re = _RAND_733[31:0];
  _RAND_734 = {1{`RANDOM}};
  _T_517_im = _RAND_734[31:0];
  _RAND_735 = {1{`RANDOM}};
  _T_518_re = _RAND_735[31:0];
  _RAND_736 = {1{`RANDOM}};
  _T_518_im = _RAND_736[31:0];
  _RAND_737 = {1{`RANDOM}};
  _T_519_re = _RAND_737[31:0];
  _RAND_738 = {1{`RANDOM}};
  _T_519_im = _RAND_738[31:0];
  _RAND_739 = {1{`RANDOM}};
  _T_520_re = _RAND_739[31:0];
  _RAND_740 = {1{`RANDOM}};
  _T_520_im = _RAND_740[31:0];
  _RAND_741 = {1{`RANDOM}};
  _T_521_re = _RAND_741[31:0];
  _RAND_742 = {1{`RANDOM}};
  _T_521_im = _RAND_742[31:0];
  _RAND_743 = {1{`RANDOM}};
  _T_522_re = _RAND_743[31:0];
  _RAND_744 = {1{`RANDOM}};
  _T_522_im = _RAND_744[31:0];
  _RAND_745 = {1{`RANDOM}};
  _T_523_re = _RAND_745[31:0];
  _RAND_746 = {1{`RANDOM}};
  _T_523_im = _RAND_746[31:0];
  _RAND_747 = {1{`RANDOM}};
  _T_524_re = _RAND_747[31:0];
  _RAND_748 = {1{`RANDOM}};
  _T_524_im = _RAND_748[31:0];
  _RAND_749 = {1{`RANDOM}};
  _T_525_re = _RAND_749[31:0];
  _RAND_750 = {1{`RANDOM}};
  _T_525_im = _RAND_750[31:0];
  _RAND_751 = {1{`RANDOM}};
  _T_526_re = _RAND_751[31:0];
  _RAND_752 = {1{`RANDOM}};
  _T_526_im = _RAND_752[31:0];
  _RAND_753 = {1{`RANDOM}};
  _T_527_re = _RAND_753[31:0];
  _RAND_754 = {1{`RANDOM}};
  _T_527_im = _RAND_754[31:0];
  _RAND_755 = {1{`RANDOM}};
  _T_528_re = _RAND_755[31:0];
  _RAND_756 = {1{`RANDOM}};
  _T_528_im = _RAND_756[31:0];
  _RAND_757 = {1{`RANDOM}};
  _T_529_re = _RAND_757[31:0];
  _RAND_758 = {1{`RANDOM}};
  _T_529_im = _RAND_758[31:0];
  _RAND_759 = {1{`RANDOM}};
  _T_530_re = _RAND_759[31:0];
  _RAND_760 = {1{`RANDOM}};
  _T_530_im = _RAND_760[31:0];
  _RAND_761 = {1{`RANDOM}};
  _T_531_re = _RAND_761[31:0];
  _RAND_762 = {1{`RANDOM}};
  _T_531_im = _RAND_762[31:0];
  _RAND_763 = {1{`RANDOM}};
  _T_532_re = _RAND_763[31:0];
  _RAND_764 = {1{`RANDOM}};
  _T_532_im = _RAND_764[31:0];
  _RAND_765 = {1{`RANDOM}};
  _T_533_re = _RAND_765[31:0];
  _RAND_766 = {1{`RANDOM}};
  _T_533_im = _RAND_766[31:0];
  _RAND_767 = {1{`RANDOM}};
  _T_534_re = _RAND_767[31:0];
  _RAND_768 = {1{`RANDOM}};
  _T_534_im = _RAND_768[31:0];
  _RAND_769 = {1{`RANDOM}};
  _T_543_re = _RAND_769[31:0];
  _RAND_770 = {1{`RANDOM}};
  _T_543_im = _RAND_770[31:0];
  _RAND_771 = {1{`RANDOM}};
  _T_544_re = _RAND_771[31:0];
  _RAND_772 = {1{`RANDOM}};
  _T_544_im = _RAND_772[31:0];
  _RAND_773 = {1{`RANDOM}};
  _T_545_re = _RAND_773[31:0];
  _RAND_774 = {1{`RANDOM}};
  _T_545_im = _RAND_774[31:0];
  _RAND_775 = {1{`RANDOM}};
  _T_546_re = _RAND_775[31:0];
  _RAND_776 = {1{`RANDOM}};
  _T_546_im = _RAND_776[31:0];
  _RAND_777 = {1{`RANDOM}};
  _T_547_re = _RAND_777[31:0];
  _RAND_778 = {1{`RANDOM}};
  _T_547_im = _RAND_778[31:0];
  _RAND_779 = {1{`RANDOM}};
  _T_548_re = _RAND_779[31:0];
  _RAND_780 = {1{`RANDOM}};
  _T_548_im = _RAND_780[31:0];
  _RAND_781 = {1{`RANDOM}};
  _T_549_re = _RAND_781[31:0];
  _RAND_782 = {1{`RANDOM}};
  _T_549_im = _RAND_782[31:0];
  _RAND_783 = {1{`RANDOM}};
  _T_550_re = _RAND_783[31:0];
  _RAND_784 = {1{`RANDOM}};
  _T_550_im = _RAND_784[31:0];
  _RAND_785 = {1{`RANDOM}};
  _T_551_re = _RAND_785[31:0];
  _RAND_786 = {1{`RANDOM}};
  _T_551_im = _RAND_786[31:0];
  _RAND_787 = {1{`RANDOM}};
  _T_552_re = _RAND_787[31:0];
  _RAND_788 = {1{`RANDOM}};
  _T_552_im = _RAND_788[31:0];
  _RAND_789 = {1{`RANDOM}};
  _T_553_re = _RAND_789[31:0];
  _RAND_790 = {1{`RANDOM}};
  _T_553_im = _RAND_790[31:0];
  _RAND_791 = {1{`RANDOM}};
  _T_554_re = _RAND_791[31:0];
  _RAND_792 = {1{`RANDOM}};
  _T_554_im = _RAND_792[31:0];
  _RAND_793 = {1{`RANDOM}};
  _T_555_re = _RAND_793[31:0];
  _RAND_794 = {1{`RANDOM}};
  _T_555_im = _RAND_794[31:0];
  _RAND_795 = {1{`RANDOM}};
  _T_556_re = _RAND_795[31:0];
  _RAND_796 = {1{`RANDOM}};
  _T_556_im = _RAND_796[31:0];
  _RAND_797 = {1{`RANDOM}};
  _T_557_re = _RAND_797[31:0];
  _RAND_798 = {1{`RANDOM}};
  _T_557_im = _RAND_798[31:0];
  _RAND_799 = {1{`RANDOM}};
  _T_558_re = _RAND_799[31:0];
  _RAND_800 = {1{`RANDOM}};
  _T_558_im = _RAND_800[31:0];
  _RAND_801 = {1{`RANDOM}};
  _T_559_re = _RAND_801[31:0];
  _RAND_802 = {1{`RANDOM}};
  _T_559_im = _RAND_802[31:0];
  _RAND_803 = {1{`RANDOM}};
  _T_560_re = _RAND_803[31:0];
  _RAND_804 = {1{`RANDOM}};
  _T_560_im = _RAND_804[31:0];
  _RAND_805 = {1{`RANDOM}};
  _T_561_re = _RAND_805[31:0];
  _RAND_806 = {1{`RANDOM}};
  _T_561_im = _RAND_806[31:0];
  _RAND_807 = {1{`RANDOM}};
  _T_562_re = _RAND_807[31:0];
  _RAND_808 = {1{`RANDOM}};
  _T_562_im = _RAND_808[31:0];
  _RAND_809 = {1{`RANDOM}};
  _T_563_re = _RAND_809[31:0];
  _RAND_810 = {1{`RANDOM}};
  _T_563_im = _RAND_810[31:0];
  _RAND_811 = {1{`RANDOM}};
  _T_564_re = _RAND_811[31:0];
  _RAND_812 = {1{`RANDOM}};
  _T_564_im = _RAND_812[31:0];
  _RAND_813 = {1{`RANDOM}};
  _T_565_re = _RAND_813[31:0];
  _RAND_814 = {1{`RANDOM}};
  _T_565_im = _RAND_814[31:0];
  _RAND_815 = {1{`RANDOM}};
  _T_566_re = _RAND_815[31:0];
  _RAND_816 = {1{`RANDOM}};
  _T_566_im = _RAND_816[31:0];
  _RAND_817 = {1{`RANDOM}};
  _T_567_re = _RAND_817[31:0];
  _RAND_818 = {1{`RANDOM}};
  _T_567_im = _RAND_818[31:0];
  _RAND_819 = {1{`RANDOM}};
  _T_568_re = _RAND_819[31:0];
  _RAND_820 = {1{`RANDOM}};
  _T_568_im = _RAND_820[31:0];
  _RAND_821 = {1{`RANDOM}};
  _T_569_re = _RAND_821[31:0];
  _RAND_822 = {1{`RANDOM}};
  _T_569_im = _RAND_822[31:0];
  _RAND_823 = {1{`RANDOM}};
  _T_570_re = _RAND_823[31:0];
  _RAND_824 = {1{`RANDOM}};
  _T_570_im = _RAND_824[31:0];
  _RAND_825 = {1{`RANDOM}};
  _T_571_re = _RAND_825[31:0];
  _RAND_826 = {1{`RANDOM}};
  _T_571_im = _RAND_826[31:0];
  _RAND_827 = {1{`RANDOM}};
  _T_572_re = _RAND_827[31:0];
  _RAND_828 = {1{`RANDOM}};
  _T_572_im = _RAND_828[31:0];
  _RAND_829 = {1{`RANDOM}};
  _T_573_re = _RAND_829[31:0];
  _RAND_830 = {1{`RANDOM}};
  _T_573_im = _RAND_830[31:0];
  _RAND_831 = {1{`RANDOM}};
  _T_574_re = _RAND_831[31:0];
  _RAND_832 = {1{`RANDOM}};
  _T_574_im = _RAND_832[31:0];
  _RAND_833 = {1{`RANDOM}};
  _T_575_re = _RAND_833[31:0];
  _RAND_834 = {1{`RANDOM}};
  _T_575_im = _RAND_834[31:0];
  _RAND_835 = {1{`RANDOM}};
  _T_576_re = _RAND_835[31:0];
  _RAND_836 = {1{`RANDOM}};
  _T_576_im = _RAND_836[31:0];
  _RAND_837 = {1{`RANDOM}};
  _T_577_re = _RAND_837[31:0];
  _RAND_838 = {1{`RANDOM}};
  _T_577_im = _RAND_838[31:0];
  _RAND_839 = {1{`RANDOM}};
  _T_578_re = _RAND_839[31:0];
  _RAND_840 = {1{`RANDOM}};
  _T_578_im = _RAND_840[31:0];
  _RAND_841 = {1{`RANDOM}};
  _T_579_re = _RAND_841[31:0];
  _RAND_842 = {1{`RANDOM}};
  _T_579_im = _RAND_842[31:0];
  _RAND_843 = {1{`RANDOM}};
  _T_580_re = _RAND_843[31:0];
  _RAND_844 = {1{`RANDOM}};
  _T_580_im = _RAND_844[31:0];
  _RAND_845 = {1{`RANDOM}};
  _T_581_re = _RAND_845[31:0];
  _RAND_846 = {1{`RANDOM}};
  _T_581_im = _RAND_846[31:0];
  _RAND_847 = {1{`RANDOM}};
  _T_582_re = _RAND_847[31:0];
  _RAND_848 = {1{`RANDOM}};
  _T_582_im = _RAND_848[31:0];
  _RAND_849 = {1{`RANDOM}};
  _T_583_re = _RAND_849[31:0];
  _RAND_850 = {1{`RANDOM}};
  _T_583_im = _RAND_850[31:0];
  _RAND_851 = {1{`RANDOM}};
  _T_584_re = _RAND_851[31:0];
  _RAND_852 = {1{`RANDOM}};
  _T_584_im = _RAND_852[31:0];
  _RAND_853 = {1{`RANDOM}};
  _T_585_re = _RAND_853[31:0];
  _RAND_854 = {1{`RANDOM}};
  _T_585_im = _RAND_854[31:0];
  _RAND_855 = {1{`RANDOM}};
  _T_586_re = _RAND_855[31:0];
  _RAND_856 = {1{`RANDOM}};
  _T_586_im = _RAND_856[31:0];
  _RAND_857 = {1{`RANDOM}};
  _T_587_re = _RAND_857[31:0];
  _RAND_858 = {1{`RANDOM}};
  _T_587_im = _RAND_858[31:0];
  _RAND_859 = {1{`RANDOM}};
  _T_588_re = _RAND_859[31:0];
  _RAND_860 = {1{`RANDOM}};
  _T_588_im = _RAND_860[31:0];
  _RAND_861 = {1{`RANDOM}};
  _T_589_re = _RAND_861[31:0];
  _RAND_862 = {1{`RANDOM}};
  _T_589_im = _RAND_862[31:0];
  _RAND_863 = {1{`RANDOM}};
  _T_590_re = _RAND_863[31:0];
  _RAND_864 = {1{`RANDOM}};
  _T_590_im = _RAND_864[31:0];
  _RAND_865 = {1{`RANDOM}};
  _T_591_re = _RAND_865[31:0];
  _RAND_866 = {1{`RANDOM}};
  _T_591_im = _RAND_866[31:0];
  _RAND_867 = {1{`RANDOM}};
  _T_592_re = _RAND_867[31:0];
  _RAND_868 = {1{`RANDOM}};
  _T_592_im = _RAND_868[31:0];
  _RAND_869 = {1{`RANDOM}};
  _T_593_re = _RAND_869[31:0];
  _RAND_870 = {1{`RANDOM}};
  _T_593_im = _RAND_870[31:0];
  _RAND_871 = {1{`RANDOM}};
  _T_594_re = _RAND_871[31:0];
  _RAND_872 = {1{`RANDOM}};
  _T_594_im = _RAND_872[31:0];
  _RAND_873 = {1{`RANDOM}};
  _T_595_re = _RAND_873[31:0];
  _RAND_874 = {1{`RANDOM}};
  _T_595_im = _RAND_874[31:0];
  _RAND_875 = {1{`RANDOM}};
  _T_596_re = _RAND_875[31:0];
  _RAND_876 = {1{`RANDOM}};
  _T_596_im = _RAND_876[31:0];
  _RAND_877 = {1{`RANDOM}};
  _T_597_re = _RAND_877[31:0];
  _RAND_878 = {1{`RANDOM}};
  _T_597_im = _RAND_878[31:0];
  _RAND_879 = {1{`RANDOM}};
  _T_598_re = _RAND_879[31:0];
  _RAND_880 = {1{`RANDOM}};
  _T_598_im = _RAND_880[31:0];
  _RAND_881 = {1{`RANDOM}};
  _T_599_re = _RAND_881[31:0];
  _RAND_882 = {1{`RANDOM}};
  _T_599_im = _RAND_882[31:0];
  _RAND_883 = {1{`RANDOM}};
  _T_600_re = _RAND_883[31:0];
  _RAND_884 = {1{`RANDOM}};
  _T_600_im = _RAND_884[31:0];
  _RAND_885 = {1{`RANDOM}};
  _T_601_re = _RAND_885[31:0];
  _RAND_886 = {1{`RANDOM}};
  _T_601_im = _RAND_886[31:0];
  _RAND_887 = {1{`RANDOM}};
  _T_602_re = _RAND_887[31:0];
  _RAND_888 = {1{`RANDOM}};
  _T_602_im = _RAND_888[31:0];
  _RAND_889 = {1{`RANDOM}};
  _T_603_re = _RAND_889[31:0];
  _RAND_890 = {1{`RANDOM}};
  _T_603_im = _RAND_890[31:0];
  _RAND_891 = {1{`RANDOM}};
  _T_604_re = _RAND_891[31:0];
  _RAND_892 = {1{`RANDOM}};
  _T_604_im = _RAND_892[31:0];
  _RAND_893 = {1{`RANDOM}};
  _T_605_re = _RAND_893[31:0];
  _RAND_894 = {1{`RANDOM}};
  _T_605_im = _RAND_894[31:0];
  _RAND_895 = {1{`RANDOM}};
  _T_606_re = _RAND_895[31:0];
  _RAND_896 = {1{`RANDOM}};
  _T_606_im = _RAND_896[31:0];
  _RAND_897 = {1{`RANDOM}};
  _T_607_re = _RAND_897[31:0];
  _RAND_898 = {1{`RANDOM}};
  _T_607_im = _RAND_898[31:0];
  _RAND_899 = {1{`RANDOM}};
  _T_608_re = _RAND_899[31:0];
  _RAND_900 = {1{`RANDOM}};
  _T_608_im = _RAND_900[31:0];
  _RAND_901 = {1{`RANDOM}};
  _T_609_re = _RAND_901[31:0];
  _RAND_902 = {1{`RANDOM}};
  _T_609_im = _RAND_902[31:0];
  _RAND_903 = {1{`RANDOM}};
  _T_610_re = _RAND_903[31:0];
  _RAND_904 = {1{`RANDOM}};
  _T_610_im = _RAND_904[31:0];
  _RAND_905 = {1{`RANDOM}};
  _T_611_re = _RAND_905[31:0];
  _RAND_906 = {1{`RANDOM}};
  _T_611_im = _RAND_906[31:0];
  _RAND_907 = {1{`RANDOM}};
  _T_612_re = _RAND_907[31:0];
  _RAND_908 = {1{`RANDOM}};
  _T_612_im = _RAND_908[31:0];
  _RAND_909 = {1{`RANDOM}};
  _T_613_re = _RAND_909[31:0];
  _RAND_910 = {1{`RANDOM}};
  _T_613_im = _RAND_910[31:0];
  _RAND_911 = {1{`RANDOM}};
  _T_614_re = _RAND_911[31:0];
  _RAND_912 = {1{`RANDOM}};
  _T_614_im = _RAND_912[31:0];
  _RAND_913 = {1{`RANDOM}};
  _T_615_re = _RAND_913[31:0];
  _RAND_914 = {1{`RANDOM}};
  _T_615_im = _RAND_914[31:0];
  _RAND_915 = {1{`RANDOM}};
  _T_616_re = _RAND_915[31:0];
  _RAND_916 = {1{`RANDOM}};
  _T_616_im = _RAND_916[31:0];
  _RAND_917 = {1{`RANDOM}};
  _T_617_re = _RAND_917[31:0];
  _RAND_918 = {1{`RANDOM}};
  _T_617_im = _RAND_918[31:0];
  _RAND_919 = {1{`RANDOM}};
  _T_618_re = _RAND_919[31:0];
  _RAND_920 = {1{`RANDOM}};
  _T_618_im = _RAND_920[31:0];
  _RAND_921 = {1{`RANDOM}};
  _T_619_re = _RAND_921[31:0];
  _RAND_922 = {1{`RANDOM}};
  _T_619_im = _RAND_922[31:0];
  _RAND_923 = {1{`RANDOM}};
  _T_620_re = _RAND_923[31:0];
  _RAND_924 = {1{`RANDOM}};
  _T_620_im = _RAND_924[31:0];
  _RAND_925 = {1{`RANDOM}};
  _T_621_re = _RAND_925[31:0];
  _RAND_926 = {1{`RANDOM}};
  _T_621_im = _RAND_926[31:0];
  _RAND_927 = {1{`RANDOM}};
  _T_622_re = _RAND_927[31:0];
  _RAND_928 = {1{`RANDOM}};
  _T_622_im = _RAND_928[31:0];
  _RAND_929 = {1{`RANDOM}};
  _T_623_re = _RAND_929[31:0];
  _RAND_930 = {1{`RANDOM}};
  _T_623_im = _RAND_930[31:0];
  _RAND_931 = {1{`RANDOM}};
  _T_624_re = _RAND_931[31:0];
  _RAND_932 = {1{`RANDOM}};
  _T_624_im = _RAND_932[31:0];
  _RAND_933 = {1{`RANDOM}};
  _T_625_re = _RAND_933[31:0];
  _RAND_934 = {1{`RANDOM}};
  _T_625_im = _RAND_934[31:0];
  _RAND_935 = {1{`RANDOM}};
  _T_626_re = _RAND_935[31:0];
  _RAND_936 = {1{`RANDOM}};
  _T_626_im = _RAND_936[31:0];
  _RAND_937 = {1{`RANDOM}};
  _T_627_re = _RAND_937[31:0];
  _RAND_938 = {1{`RANDOM}};
  _T_627_im = _RAND_938[31:0];
  _RAND_939 = {1{`RANDOM}};
  _T_628_re = _RAND_939[31:0];
  _RAND_940 = {1{`RANDOM}};
  _T_628_im = _RAND_940[31:0];
  _RAND_941 = {1{`RANDOM}};
  _T_629_re = _RAND_941[31:0];
  _RAND_942 = {1{`RANDOM}};
  _T_629_im = _RAND_942[31:0];
  _RAND_943 = {1{`RANDOM}};
  _T_630_re = _RAND_943[31:0];
  _RAND_944 = {1{`RANDOM}};
  _T_630_im = _RAND_944[31:0];
  _RAND_945 = {1{`RANDOM}};
  _T_631_re = _RAND_945[31:0];
  _RAND_946 = {1{`RANDOM}};
  _T_631_im = _RAND_946[31:0];
  _RAND_947 = {1{`RANDOM}};
  _T_632_re = _RAND_947[31:0];
  _RAND_948 = {1{`RANDOM}};
  _T_632_im = _RAND_948[31:0];
  _RAND_949 = {1{`RANDOM}};
  _T_633_re = _RAND_949[31:0];
  _RAND_950 = {1{`RANDOM}};
  _T_633_im = _RAND_950[31:0];
  _RAND_951 = {1{`RANDOM}};
  _T_634_re = _RAND_951[31:0];
  _RAND_952 = {1{`RANDOM}};
  _T_634_im = _RAND_952[31:0];
  _RAND_953 = {1{`RANDOM}};
  _T_635_re = _RAND_953[31:0];
  _RAND_954 = {1{`RANDOM}};
  _T_635_im = _RAND_954[31:0];
  _RAND_955 = {1{`RANDOM}};
  _T_636_re = _RAND_955[31:0];
  _RAND_956 = {1{`RANDOM}};
  _T_636_im = _RAND_956[31:0];
  _RAND_957 = {1{`RANDOM}};
  _T_637_re = _RAND_957[31:0];
  _RAND_958 = {1{`RANDOM}};
  _T_637_im = _RAND_958[31:0];
  _RAND_959 = {1{`RANDOM}};
  _T_638_re = _RAND_959[31:0];
  _RAND_960 = {1{`RANDOM}};
  _T_638_im = _RAND_960[31:0];
  _RAND_961 = {1{`RANDOM}};
  _T_639_re = _RAND_961[31:0];
  _RAND_962 = {1{`RANDOM}};
  _T_639_im = _RAND_962[31:0];
  _RAND_963 = {1{`RANDOM}};
  _T_640_re = _RAND_963[31:0];
  _RAND_964 = {1{`RANDOM}};
  _T_640_im = _RAND_964[31:0];
  _RAND_965 = {1{`RANDOM}};
  _T_641_re = _RAND_965[31:0];
  _RAND_966 = {1{`RANDOM}};
  _T_641_im = _RAND_966[31:0];
  _RAND_967 = {1{`RANDOM}};
  _T_642_re = _RAND_967[31:0];
  _RAND_968 = {1{`RANDOM}};
  _T_642_im = _RAND_968[31:0];
  _RAND_969 = {1{`RANDOM}};
  _T_643_re = _RAND_969[31:0];
  _RAND_970 = {1{`RANDOM}};
  _T_643_im = _RAND_970[31:0];
  _RAND_971 = {1{`RANDOM}};
  _T_644_re = _RAND_971[31:0];
  _RAND_972 = {1{`RANDOM}};
  _T_644_im = _RAND_972[31:0];
  _RAND_973 = {1{`RANDOM}};
  _T_645_re = _RAND_973[31:0];
  _RAND_974 = {1{`RANDOM}};
  _T_645_im = _RAND_974[31:0];
  _RAND_975 = {1{`RANDOM}};
  _T_646_re = _RAND_975[31:0];
  _RAND_976 = {1{`RANDOM}};
  _T_646_im = _RAND_976[31:0];
  _RAND_977 = {1{`RANDOM}};
  _T_647_re = _RAND_977[31:0];
  _RAND_978 = {1{`RANDOM}};
  _T_647_im = _RAND_978[31:0];
  _RAND_979 = {1{`RANDOM}};
  _T_648_re = _RAND_979[31:0];
  _RAND_980 = {1{`RANDOM}};
  _T_648_im = _RAND_980[31:0];
  _RAND_981 = {1{`RANDOM}};
  _T_649_re = _RAND_981[31:0];
  _RAND_982 = {1{`RANDOM}};
  _T_649_im = _RAND_982[31:0];
  _RAND_983 = {1{`RANDOM}};
  _T_650_re = _RAND_983[31:0];
  _RAND_984 = {1{`RANDOM}};
  _T_650_im = _RAND_984[31:0];
  _RAND_985 = {1{`RANDOM}};
  _T_651_re = _RAND_985[31:0];
  _RAND_986 = {1{`RANDOM}};
  _T_651_im = _RAND_986[31:0];
  _RAND_987 = {1{`RANDOM}};
  _T_652_re = _RAND_987[31:0];
  _RAND_988 = {1{`RANDOM}};
  _T_652_im = _RAND_988[31:0];
  _RAND_989 = {1{`RANDOM}};
  _T_653_re = _RAND_989[31:0];
  _RAND_990 = {1{`RANDOM}};
  _T_653_im = _RAND_990[31:0];
  _RAND_991 = {1{`RANDOM}};
  _T_654_re = _RAND_991[31:0];
  _RAND_992 = {1{`RANDOM}};
  _T_654_im = _RAND_992[31:0];
  _RAND_993 = {1{`RANDOM}};
  _T_655_re = _RAND_993[31:0];
  _RAND_994 = {1{`RANDOM}};
  _T_655_im = _RAND_994[31:0];
  _RAND_995 = {1{`RANDOM}};
  _T_656_re = _RAND_995[31:0];
  _RAND_996 = {1{`RANDOM}};
  _T_656_im = _RAND_996[31:0];
  _RAND_997 = {1{`RANDOM}};
  _T_657_re = _RAND_997[31:0];
  _RAND_998 = {1{`RANDOM}};
  _T_657_im = _RAND_998[31:0];
  _RAND_999 = {1{`RANDOM}};
  _T_658_re = _RAND_999[31:0];
  _RAND_1000 = {1{`RANDOM}};
  _T_658_im = _RAND_1000[31:0];
  _RAND_1001 = {1{`RANDOM}};
  _T_659_re = _RAND_1001[31:0];
  _RAND_1002 = {1{`RANDOM}};
  _T_659_im = _RAND_1002[31:0];
  _RAND_1003 = {1{`RANDOM}};
  _T_660_re = _RAND_1003[31:0];
  _RAND_1004 = {1{`RANDOM}};
  _T_660_im = _RAND_1004[31:0];
  _RAND_1005 = {1{`RANDOM}};
  _T_661_re = _RAND_1005[31:0];
  _RAND_1006 = {1{`RANDOM}};
  _T_661_im = _RAND_1006[31:0];
  _RAND_1007 = {1{`RANDOM}};
  _T_662_re = _RAND_1007[31:0];
  _RAND_1008 = {1{`RANDOM}};
  _T_662_im = _RAND_1008[31:0];
  _RAND_1009 = {1{`RANDOM}};
  _T_663_re = _RAND_1009[31:0];
  _RAND_1010 = {1{`RANDOM}};
  _T_663_im = _RAND_1010[31:0];
  _RAND_1011 = {1{`RANDOM}};
  _T_664_re = _RAND_1011[31:0];
  _RAND_1012 = {1{`RANDOM}};
  _T_664_im = _RAND_1012[31:0];
  _RAND_1013 = {1{`RANDOM}};
  _T_665_re = _RAND_1013[31:0];
  _RAND_1014 = {1{`RANDOM}};
  _T_665_im = _RAND_1014[31:0];
  _RAND_1015 = {1{`RANDOM}};
  _T_666_re = _RAND_1015[31:0];
  _RAND_1016 = {1{`RANDOM}};
  _T_666_im = _RAND_1016[31:0];
  _RAND_1017 = {1{`RANDOM}};
  _T_667_re = _RAND_1017[31:0];
  _RAND_1018 = {1{`RANDOM}};
  _T_667_im = _RAND_1018[31:0];
  _RAND_1019 = {1{`RANDOM}};
  _T_668_re = _RAND_1019[31:0];
  _RAND_1020 = {1{`RANDOM}};
  _T_668_im = _RAND_1020[31:0];
  _RAND_1021 = {1{`RANDOM}};
  _T_669_re = _RAND_1021[31:0];
  _RAND_1022 = {1{`RANDOM}};
  _T_669_im = _RAND_1022[31:0];
  _RAND_1023 = {1{`RANDOM}};
  _T_670_re = _RAND_1023[31:0];
  _RAND_1024 = {1{`RANDOM}};
  _T_670_im = _RAND_1024[31:0];
  _RAND_1025 = {1{`RANDOM}};
  _T_672_re = _RAND_1025[31:0];
  _RAND_1026 = {1{`RANDOM}};
  _T_672_im = _RAND_1026[31:0];
  _RAND_1027 = {1{`RANDOM}};
  _T_673_re = _RAND_1027[31:0];
  _RAND_1028 = {1{`RANDOM}};
  _T_673_im = _RAND_1028[31:0];
  _RAND_1029 = {1{`RANDOM}};
  _T_674_re = _RAND_1029[31:0];
  _RAND_1030 = {1{`RANDOM}};
  _T_674_im = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  _T_675_re = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  _T_675_im = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  _T_676_re = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  _T_676_im = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  _T_677_re = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  _T_677_im = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  _T_678_re = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  _T_678_im = _RAND_1038[31:0];
  _RAND_1039 = {1{`RANDOM}};
  _T_679_re = _RAND_1039[31:0];
  _RAND_1040 = {1{`RANDOM}};
  _T_679_im = _RAND_1040[31:0];
  _RAND_1041 = {1{`RANDOM}};
  _T_680_re = _RAND_1041[31:0];
  _RAND_1042 = {1{`RANDOM}};
  _T_680_im = _RAND_1042[31:0];
  _RAND_1043 = {1{`RANDOM}};
  _T_681_re = _RAND_1043[31:0];
  _RAND_1044 = {1{`RANDOM}};
  _T_681_im = _RAND_1044[31:0];
  _RAND_1045 = {1{`RANDOM}};
  _T_682_re = _RAND_1045[31:0];
  _RAND_1046 = {1{`RANDOM}};
  _T_682_im = _RAND_1046[31:0];
  _RAND_1047 = {1{`RANDOM}};
  _T_683_re = _RAND_1047[31:0];
  _RAND_1048 = {1{`RANDOM}};
  _T_683_im = _RAND_1048[31:0];
  _RAND_1049 = {1{`RANDOM}};
  _T_684_re = _RAND_1049[31:0];
  _RAND_1050 = {1{`RANDOM}};
  _T_684_im = _RAND_1050[31:0];
  _RAND_1051 = {1{`RANDOM}};
  _T_685_re = _RAND_1051[31:0];
  _RAND_1052 = {1{`RANDOM}};
  _T_685_im = _RAND_1052[31:0];
  _RAND_1053 = {1{`RANDOM}};
  _T_686_re = _RAND_1053[31:0];
  _RAND_1054 = {1{`RANDOM}};
  _T_686_im = _RAND_1054[31:0];
  _RAND_1055 = {1{`RANDOM}};
  _T_687_re = _RAND_1055[31:0];
  _RAND_1056 = {1{`RANDOM}};
  _T_687_im = _RAND_1056[31:0];
  _RAND_1057 = {1{`RANDOM}};
  _T_688_re = _RAND_1057[31:0];
  _RAND_1058 = {1{`RANDOM}};
  _T_688_im = _RAND_1058[31:0];
  _RAND_1059 = {1{`RANDOM}};
  _T_689_re = _RAND_1059[31:0];
  _RAND_1060 = {1{`RANDOM}};
  _T_689_im = _RAND_1060[31:0];
  _RAND_1061 = {1{`RANDOM}};
  _T_690_re = _RAND_1061[31:0];
  _RAND_1062 = {1{`RANDOM}};
  _T_690_im = _RAND_1062[31:0];
  _RAND_1063 = {1{`RANDOM}};
  _T_691_re = _RAND_1063[31:0];
  _RAND_1064 = {1{`RANDOM}};
  _T_691_im = _RAND_1064[31:0];
  _RAND_1065 = {1{`RANDOM}};
  _T_692_re = _RAND_1065[31:0];
  _RAND_1066 = {1{`RANDOM}};
  _T_692_im = _RAND_1066[31:0];
  _RAND_1067 = {1{`RANDOM}};
  _T_693_re = _RAND_1067[31:0];
  _RAND_1068 = {1{`RANDOM}};
  _T_693_im = _RAND_1068[31:0];
  _RAND_1069 = {1{`RANDOM}};
  _T_694_re = _RAND_1069[31:0];
  _RAND_1070 = {1{`RANDOM}};
  _T_694_im = _RAND_1070[31:0];
  _RAND_1071 = {1{`RANDOM}};
  _T_695_re = _RAND_1071[31:0];
  _RAND_1072 = {1{`RANDOM}};
  _T_695_im = _RAND_1072[31:0];
  _RAND_1073 = {1{`RANDOM}};
  _T_696_re = _RAND_1073[31:0];
  _RAND_1074 = {1{`RANDOM}};
  _T_696_im = _RAND_1074[31:0];
  _RAND_1075 = {1{`RANDOM}};
  _T_697_re = _RAND_1075[31:0];
  _RAND_1076 = {1{`RANDOM}};
  _T_697_im = _RAND_1076[31:0];
  _RAND_1077 = {1{`RANDOM}};
  _T_698_re = _RAND_1077[31:0];
  _RAND_1078 = {1{`RANDOM}};
  _T_698_im = _RAND_1078[31:0];
  _RAND_1079 = {1{`RANDOM}};
  _T_699_re = _RAND_1079[31:0];
  _RAND_1080 = {1{`RANDOM}};
  _T_699_im = _RAND_1080[31:0];
  _RAND_1081 = {1{`RANDOM}};
  _T_700_re = _RAND_1081[31:0];
  _RAND_1082 = {1{`RANDOM}};
  _T_700_im = _RAND_1082[31:0];
  _RAND_1083 = {1{`RANDOM}};
  _T_701_re = _RAND_1083[31:0];
  _RAND_1084 = {1{`RANDOM}};
  _T_701_im = _RAND_1084[31:0];
  _RAND_1085 = {1{`RANDOM}};
  _T_702_re = _RAND_1085[31:0];
  _RAND_1086 = {1{`RANDOM}};
  _T_702_im = _RAND_1086[31:0];
  _RAND_1087 = {1{`RANDOM}};
  _T_703_re = _RAND_1087[31:0];
  _RAND_1088 = {1{`RANDOM}};
  _T_703_im = _RAND_1088[31:0];
  _RAND_1089 = {1{`RANDOM}};
  _T_704_re = _RAND_1089[31:0];
  _RAND_1090 = {1{`RANDOM}};
  _T_704_im = _RAND_1090[31:0];
  _RAND_1091 = {1{`RANDOM}};
  _T_705_re = _RAND_1091[31:0];
  _RAND_1092 = {1{`RANDOM}};
  _T_705_im = _RAND_1092[31:0];
  _RAND_1093 = {1{`RANDOM}};
  _T_706_re = _RAND_1093[31:0];
  _RAND_1094 = {1{`RANDOM}};
  _T_706_im = _RAND_1094[31:0];
  _RAND_1095 = {1{`RANDOM}};
  _T_707_re = _RAND_1095[31:0];
  _RAND_1096 = {1{`RANDOM}};
  _T_707_im = _RAND_1096[31:0];
  _RAND_1097 = {1{`RANDOM}};
  _T_708_re = _RAND_1097[31:0];
  _RAND_1098 = {1{`RANDOM}};
  _T_708_im = _RAND_1098[31:0];
  _RAND_1099 = {1{`RANDOM}};
  _T_709_re = _RAND_1099[31:0];
  _RAND_1100 = {1{`RANDOM}};
  _T_709_im = _RAND_1100[31:0];
  _RAND_1101 = {1{`RANDOM}};
  _T_710_re = _RAND_1101[31:0];
  _RAND_1102 = {1{`RANDOM}};
  _T_710_im = _RAND_1102[31:0];
  _RAND_1103 = {1{`RANDOM}};
  _T_711_re = _RAND_1103[31:0];
  _RAND_1104 = {1{`RANDOM}};
  _T_711_im = _RAND_1104[31:0];
  _RAND_1105 = {1{`RANDOM}};
  _T_712_re = _RAND_1105[31:0];
  _RAND_1106 = {1{`RANDOM}};
  _T_712_im = _RAND_1106[31:0];
  _RAND_1107 = {1{`RANDOM}};
  _T_713_re = _RAND_1107[31:0];
  _RAND_1108 = {1{`RANDOM}};
  _T_713_im = _RAND_1108[31:0];
  _RAND_1109 = {1{`RANDOM}};
  _T_714_re = _RAND_1109[31:0];
  _RAND_1110 = {1{`RANDOM}};
  _T_714_im = _RAND_1110[31:0];
  _RAND_1111 = {1{`RANDOM}};
  _T_715_re = _RAND_1111[31:0];
  _RAND_1112 = {1{`RANDOM}};
  _T_715_im = _RAND_1112[31:0];
  _RAND_1113 = {1{`RANDOM}};
  _T_716_re = _RAND_1113[31:0];
  _RAND_1114 = {1{`RANDOM}};
  _T_716_im = _RAND_1114[31:0];
  _RAND_1115 = {1{`RANDOM}};
  _T_717_re = _RAND_1115[31:0];
  _RAND_1116 = {1{`RANDOM}};
  _T_717_im = _RAND_1116[31:0];
  _RAND_1117 = {1{`RANDOM}};
  _T_718_re = _RAND_1117[31:0];
  _RAND_1118 = {1{`RANDOM}};
  _T_718_im = _RAND_1118[31:0];
  _RAND_1119 = {1{`RANDOM}};
  _T_719_re = _RAND_1119[31:0];
  _RAND_1120 = {1{`RANDOM}};
  _T_719_im = _RAND_1120[31:0];
  _RAND_1121 = {1{`RANDOM}};
  _T_720_re = _RAND_1121[31:0];
  _RAND_1122 = {1{`RANDOM}};
  _T_720_im = _RAND_1122[31:0];
  _RAND_1123 = {1{`RANDOM}};
  _T_721_re = _RAND_1123[31:0];
  _RAND_1124 = {1{`RANDOM}};
  _T_721_im = _RAND_1124[31:0];
  _RAND_1125 = {1{`RANDOM}};
  _T_722_re = _RAND_1125[31:0];
  _RAND_1126 = {1{`RANDOM}};
  _T_722_im = _RAND_1126[31:0];
  _RAND_1127 = {1{`RANDOM}};
  _T_723_re = _RAND_1127[31:0];
  _RAND_1128 = {1{`RANDOM}};
  _T_723_im = _RAND_1128[31:0];
  _RAND_1129 = {1{`RANDOM}};
  _T_724_re = _RAND_1129[31:0];
  _RAND_1130 = {1{`RANDOM}};
  _T_724_im = _RAND_1130[31:0];
  _RAND_1131 = {1{`RANDOM}};
  _T_725_re = _RAND_1131[31:0];
  _RAND_1132 = {1{`RANDOM}};
  _T_725_im = _RAND_1132[31:0];
  _RAND_1133 = {1{`RANDOM}};
  _T_726_re = _RAND_1133[31:0];
  _RAND_1134 = {1{`RANDOM}};
  _T_726_im = _RAND_1134[31:0];
  _RAND_1135 = {1{`RANDOM}};
  _T_727_re = _RAND_1135[31:0];
  _RAND_1136 = {1{`RANDOM}};
  _T_727_im = _RAND_1136[31:0];
  _RAND_1137 = {1{`RANDOM}};
  _T_728_re = _RAND_1137[31:0];
  _RAND_1138 = {1{`RANDOM}};
  _T_728_im = _RAND_1138[31:0];
  _RAND_1139 = {1{`RANDOM}};
  _T_729_re = _RAND_1139[31:0];
  _RAND_1140 = {1{`RANDOM}};
  _T_729_im = _RAND_1140[31:0];
  _RAND_1141 = {1{`RANDOM}};
  _T_730_re = _RAND_1141[31:0];
  _RAND_1142 = {1{`RANDOM}};
  _T_730_im = _RAND_1142[31:0];
  _RAND_1143 = {1{`RANDOM}};
  _T_731_re = _RAND_1143[31:0];
  _RAND_1144 = {1{`RANDOM}};
  _T_731_im = _RAND_1144[31:0];
  _RAND_1145 = {1{`RANDOM}};
  _T_732_re = _RAND_1145[31:0];
  _RAND_1146 = {1{`RANDOM}};
  _T_732_im = _RAND_1146[31:0];
  _RAND_1147 = {1{`RANDOM}};
  _T_733_re = _RAND_1147[31:0];
  _RAND_1148 = {1{`RANDOM}};
  _T_733_im = _RAND_1148[31:0];
  _RAND_1149 = {1{`RANDOM}};
  _T_734_re = _RAND_1149[31:0];
  _RAND_1150 = {1{`RANDOM}};
  _T_734_im = _RAND_1150[31:0];
  _RAND_1151 = {1{`RANDOM}};
  _T_735_re = _RAND_1151[31:0];
  _RAND_1152 = {1{`RANDOM}};
  _T_735_im = _RAND_1152[31:0];
  _RAND_1153 = {1{`RANDOM}};
  _T_744_re = _RAND_1153[31:0];
  _RAND_1154 = {1{`RANDOM}};
  _T_744_im = _RAND_1154[31:0];
  _RAND_1155 = {1{`RANDOM}};
  _T_745_re = _RAND_1155[31:0];
  _RAND_1156 = {1{`RANDOM}};
  _T_745_im = _RAND_1156[31:0];
  _RAND_1157 = {1{`RANDOM}};
  _T_746_re = _RAND_1157[31:0];
  _RAND_1158 = {1{`RANDOM}};
  _T_746_im = _RAND_1158[31:0];
  _RAND_1159 = {1{`RANDOM}};
  _T_747_re = _RAND_1159[31:0];
  _RAND_1160 = {1{`RANDOM}};
  _T_747_im = _RAND_1160[31:0];
  _RAND_1161 = {1{`RANDOM}};
  _T_748_re = _RAND_1161[31:0];
  _RAND_1162 = {1{`RANDOM}};
  _T_748_im = _RAND_1162[31:0];
  _RAND_1163 = {1{`RANDOM}};
  _T_749_re = _RAND_1163[31:0];
  _RAND_1164 = {1{`RANDOM}};
  _T_749_im = _RAND_1164[31:0];
  _RAND_1165 = {1{`RANDOM}};
  _T_750_re = _RAND_1165[31:0];
  _RAND_1166 = {1{`RANDOM}};
  _T_750_im = _RAND_1166[31:0];
  _RAND_1167 = {1{`RANDOM}};
  _T_751_re = _RAND_1167[31:0];
  _RAND_1168 = {1{`RANDOM}};
  _T_751_im = _RAND_1168[31:0];
  _RAND_1169 = {1{`RANDOM}};
  _T_752_re = _RAND_1169[31:0];
  _RAND_1170 = {1{`RANDOM}};
  _T_752_im = _RAND_1170[31:0];
  _RAND_1171 = {1{`RANDOM}};
  _T_753_re = _RAND_1171[31:0];
  _RAND_1172 = {1{`RANDOM}};
  _T_753_im = _RAND_1172[31:0];
  _RAND_1173 = {1{`RANDOM}};
  _T_754_re = _RAND_1173[31:0];
  _RAND_1174 = {1{`RANDOM}};
  _T_754_im = _RAND_1174[31:0];
  _RAND_1175 = {1{`RANDOM}};
  _T_755_re = _RAND_1175[31:0];
  _RAND_1176 = {1{`RANDOM}};
  _T_755_im = _RAND_1176[31:0];
  _RAND_1177 = {1{`RANDOM}};
  _T_756_re = _RAND_1177[31:0];
  _RAND_1178 = {1{`RANDOM}};
  _T_756_im = _RAND_1178[31:0];
  _RAND_1179 = {1{`RANDOM}};
  _T_757_re = _RAND_1179[31:0];
  _RAND_1180 = {1{`RANDOM}};
  _T_757_im = _RAND_1180[31:0];
  _RAND_1181 = {1{`RANDOM}};
  _T_758_re = _RAND_1181[31:0];
  _RAND_1182 = {1{`RANDOM}};
  _T_758_im = _RAND_1182[31:0];
  _RAND_1183 = {1{`RANDOM}};
  _T_759_re = _RAND_1183[31:0];
  _RAND_1184 = {1{`RANDOM}};
  _T_759_im = _RAND_1184[31:0];
  _RAND_1185 = {1{`RANDOM}};
  _T_760_re = _RAND_1185[31:0];
  _RAND_1186 = {1{`RANDOM}};
  _T_760_im = _RAND_1186[31:0];
  _RAND_1187 = {1{`RANDOM}};
  _T_761_re = _RAND_1187[31:0];
  _RAND_1188 = {1{`RANDOM}};
  _T_761_im = _RAND_1188[31:0];
  _RAND_1189 = {1{`RANDOM}};
  _T_762_re = _RAND_1189[31:0];
  _RAND_1190 = {1{`RANDOM}};
  _T_762_im = _RAND_1190[31:0];
  _RAND_1191 = {1{`RANDOM}};
  _T_763_re = _RAND_1191[31:0];
  _RAND_1192 = {1{`RANDOM}};
  _T_763_im = _RAND_1192[31:0];
  _RAND_1193 = {1{`RANDOM}};
  _T_764_re = _RAND_1193[31:0];
  _RAND_1194 = {1{`RANDOM}};
  _T_764_im = _RAND_1194[31:0];
  _RAND_1195 = {1{`RANDOM}};
  _T_765_re = _RAND_1195[31:0];
  _RAND_1196 = {1{`RANDOM}};
  _T_765_im = _RAND_1196[31:0];
  _RAND_1197 = {1{`RANDOM}};
  _T_766_re = _RAND_1197[31:0];
  _RAND_1198 = {1{`RANDOM}};
  _T_766_im = _RAND_1198[31:0];
  _RAND_1199 = {1{`RANDOM}};
  _T_767_re = _RAND_1199[31:0];
  _RAND_1200 = {1{`RANDOM}};
  _T_767_im = _RAND_1200[31:0];
  _RAND_1201 = {1{`RANDOM}};
  _T_768_re = _RAND_1201[31:0];
  _RAND_1202 = {1{`RANDOM}};
  _T_768_im = _RAND_1202[31:0];
  _RAND_1203 = {1{`RANDOM}};
  _T_769_re = _RAND_1203[31:0];
  _RAND_1204 = {1{`RANDOM}};
  _T_769_im = _RAND_1204[31:0];
  _RAND_1205 = {1{`RANDOM}};
  _T_770_re = _RAND_1205[31:0];
  _RAND_1206 = {1{`RANDOM}};
  _T_770_im = _RAND_1206[31:0];
  _RAND_1207 = {1{`RANDOM}};
  _T_771_re = _RAND_1207[31:0];
  _RAND_1208 = {1{`RANDOM}};
  _T_771_im = _RAND_1208[31:0];
  _RAND_1209 = {1{`RANDOM}};
  _T_772_re = _RAND_1209[31:0];
  _RAND_1210 = {1{`RANDOM}};
  _T_772_im = _RAND_1210[31:0];
  _RAND_1211 = {1{`RANDOM}};
  _T_773_re = _RAND_1211[31:0];
  _RAND_1212 = {1{`RANDOM}};
  _T_773_im = _RAND_1212[31:0];
  _RAND_1213 = {1{`RANDOM}};
  _T_774_re = _RAND_1213[31:0];
  _RAND_1214 = {1{`RANDOM}};
  _T_774_im = _RAND_1214[31:0];
  _RAND_1215 = {1{`RANDOM}};
  _T_775_re = _RAND_1215[31:0];
  _RAND_1216 = {1{`RANDOM}};
  _T_775_im = _RAND_1216[31:0];
  _RAND_1217 = {1{`RANDOM}};
  _T_776_re = _RAND_1217[31:0];
  _RAND_1218 = {1{`RANDOM}};
  _T_776_im = _RAND_1218[31:0];
  _RAND_1219 = {1{`RANDOM}};
  _T_777_re = _RAND_1219[31:0];
  _RAND_1220 = {1{`RANDOM}};
  _T_777_im = _RAND_1220[31:0];
  _RAND_1221 = {1{`RANDOM}};
  _T_778_re = _RAND_1221[31:0];
  _RAND_1222 = {1{`RANDOM}};
  _T_778_im = _RAND_1222[31:0];
  _RAND_1223 = {1{`RANDOM}};
  _T_779_re = _RAND_1223[31:0];
  _RAND_1224 = {1{`RANDOM}};
  _T_779_im = _RAND_1224[31:0];
  _RAND_1225 = {1{`RANDOM}};
  _T_780_re = _RAND_1225[31:0];
  _RAND_1226 = {1{`RANDOM}};
  _T_780_im = _RAND_1226[31:0];
  _RAND_1227 = {1{`RANDOM}};
  _T_781_re = _RAND_1227[31:0];
  _RAND_1228 = {1{`RANDOM}};
  _T_781_im = _RAND_1228[31:0];
  _RAND_1229 = {1{`RANDOM}};
  _T_782_re = _RAND_1229[31:0];
  _RAND_1230 = {1{`RANDOM}};
  _T_782_im = _RAND_1230[31:0];
  _RAND_1231 = {1{`RANDOM}};
  _T_783_re = _RAND_1231[31:0];
  _RAND_1232 = {1{`RANDOM}};
  _T_783_im = _RAND_1232[31:0];
  _RAND_1233 = {1{`RANDOM}};
  _T_784_re = _RAND_1233[31:0];
  _RAND_1234 = {1{`RANDOM}};
  _T_784_im = _RAND_1234[31:0];
  _RAND_1235 = {1{`RANDOM}};
  _T_785_re = _RAND_1235[31:0];
  _RAND_1236 = {1{`RANDOM}};
  _T_785_im = _RAND_1236[31:0];
  _RAND_1237 = {1{`RANDOM}};
  _T_786_re = _RAND_1237[31:0];
  _RAND_1238 = {1{`RANDOM}};
  _T_786_im = _RAND_1238[31:0];
  _RAND_1239 = {1{`RANDOM}};
  _T_787_re = _RAND_1239[31:0];
  _RAND_1240 = {1{`RANDOM}};
  _T_787_im = _RAND_1240[31:0];
  _RAND_1241 = {1{`RANDOM}};
  _T_788_re = _RAND_1241[31:0];
  _RAND_1242 = {1{`RANDOM}};
  _T_788_im = _RAND_1242[31:0];
  _RAND_1243 = {1{`RANDOM}};
  _T_789_re = _RAND_1243[31:0];
  _RAND_1244 = {1{`RANDOM}};
  _T_789_im = _RAND_1244[31:0];
  _RAND_1245 = {1{`RANDOM}};
  _T_790_re = _RAND_1245[31:0];
  _RAND_1246 = {1{`RANDOM}};
  _T_790_im = _RAND_1246[31:0];
  _RAND_1247 = {1{`RANDOM}};
  _T_791_re = _RAND_1247[31:0];
  _RAND_1248 = {1{`RANDOM}};
  _T_791_im = _RAND_1248[31:0];
  _RAND_1249 = {1{`RANDOM}};
  _T_792_re = _RAND_1249[31:0];
  _RAND_1250 = {1{`RANDOM}};
  _T_792_im = _RAND_1250[31:0];
  _RAND_1251 = {1{`RANDOM}};
  _T_793_re = _RAND_1251[31:0];
  _RAND_1252 = {1{`RANDOM}};
  _T_793_im = _RAND_1252[31:0];
  _RAND_1253 = {1{`RANDOM}};
  _T_794_re = _RAND_1253[31:0];
  _RAND_1254 = {1{`RANDOM}};
  _T_794_im = _RAND_1254[31:0];
  _RAND_1255 = {1{`RANDOM}};
  _T_795_re = _RAND_1255[31:0];
  _RAND_1256 = {1{`RANDOM}};
  _T_795_im = _RAND_1256[31:0];
  _RAND_1257 = {1{`RANDOM}};
  _T_796_re = _RAND_1257[31:0];
  _RAND_1258 = {1{`RANDOM}};
  _T_796_im = _RAND_1258[31:0];
  _RAND_1259 = {1{`RANDOM}};
  _T_797_re = _RAND_1259[31:0];
  _RAND_1260 = {1{`RANDOM}};
  _T_797_im = _RAND_1260[31:0];
  _RAND_1261 = {1{`RANDOM}};
  _T_798_re = _RAND_1261[31:0];
  _RAND_1262 = {1{`RANDOM}};
  _T_798_im = _RAND_1262[31:0];
  _RAND_1263 = {1{`RANDOM}};
  _T_799_re = _RAND_1263[31:0];
  _RAND_1264 = {1{`RANDOM}};
  _T_799_im = _RAND_1264[31:0];
  _RAND_1265 = {1{`RANDOM}};
  _T_800_re = _RAND_1265[31:0];
  _RAND_1266 = {1{`RANDOM}};
  _T_800_im = _RAND_1266[31:0];
  _RAND_1267 = {1{`RANDOM}};
  _T_801_re = _RAND_1267[31:0];
  _RAND_1268 = {1{`RANDOM}};
  _T_801_im = _RAND_1268[31:0];
  _RAND_1269 = {1{`RANDOM}};
  _T_802_re = _RAND_1269[31:0];
  _RAND_1270 = {1{`RANDOM}};
  _T_802_im = _RAND_1270[31:0];
  _RAND_1271 = {1{`RANDOM}};
  _T_803_re = _RAND_1271[31:0];
  _RAND_1272 = {1{`RANDOM}};
  _T_803_im = _RAND_1272[31:0];
  _RAND_1273 = {1{`RANDOM}};
  _T_804_re = _RAND_1273[31:0];
  _RAND_1274 = {1{`RANDOM}};
  _T_804_im = _RAND_1274[31:0];
  _RAND_1275 = {1{`RANDOM}};
  _T_805_re = _RAND_1275[31:0];
  _RAND_1276 = {1{`RANDOM}};
  _T_805_im = _RAND_1276[31:0];
  _RAND_1277 = {1{`RANDOM}};
  _T_806_re = _RAND_1277[31:0];
  _RAND_1278 = {1{`RANDOM}};
  _T_806_im = _RAND_1278[31:0];
  _RAND_1279 = {1{`RANDOM}};
  _T_807_re = _RAND_1279[31:0];
  _RAND_1280 = {1{`RANDOM}};
  _T_807_im = _RAND_1280[31:0];
  _RAND_1281 = {1{`RANDOM}};
  _T_809_re = _RAND_1281[31:0];
  _RAND_1282 = {1{`RANDOM}};
  _T_809_im = _RAND_1282[31:0];
  _RAND_1283 = {1{`RANDOM}};
  _T_810_re = _RAND_1283[31:0];
  _RAND_1284 = {1{`RANDOM}};
  _T_810_im = _RAND_1284[31:0];
  _RAND_1285 = {1{`RANDOM}};
  _T_811_re = _RAND_1285[31:0];
  _RAND_1286 = {1{`RANDOM}};
  _T_811_im = _RAND_1286[31:0];
  _RAND_1287 = {1{`RANDOM}};
  _T_812_re = _RAND_1287[31:0];
  _RAND_1288 = {1{`RANDOM}};
  _T_812_im = _RAND_1288[31:0];
  _RAND_1289 = {1{`RANDOM}};
  _T_813_re = _RAND_1289[31:0];
  _RAND_1290 = {1{`RANDOM}};
  _T_813_im = _RAND_1290[31:0];
  _RAND_1291 = {1{`RANDOM}};
  _T_814_re = _RAND_1291[31:0];
  _RAND_1292 = {1{`RANDOM}};
  _T_814_im = _RAND_1292[31:0];
  _RAND_1293 = {1{`RANDOM}};
  _T_815_re = _RAND_1293[31:0];
  _RAND_1294 = {1{`RANDOM}};
  _T_815_im = _RAND_1294[31:0];
  _RAND_1295 = {1{`RANDOM}};
  _T_816_re = _RAND_1295[31:0];
  _RAND_1296 = {1{`RANDOM}};
  _T_816_im = _RAND_1296[31:0];
  _RAND_1297 = {1{`RANDOM}};
  _T_817_re = _RAND_1297[31:0];
  _RAND_1298 = {1{`RANDOM}};
  _T_817_im = _RAND_1298[31:0];
  _RAND_1299 = {1{`RANDOM}};
  _T_818_re = _RAND_1299[31:0];
  _RAND_1300 = {1{`RANDOM}};
  _T_818_im = _RAND_1300[31:0];
  _RAND_1301 = {1{`RANDOM}};
  _T_819_re = _RAND_1301[31:0];
  _RAND_1302 = {1{`RANDOM}};
  _T_819_im = _RAND_1302[31:0];
  _RAND_1303 = {1{`RANDOM}};
  _T_820_re = _RAND_1303[31:0];
  _RAND_1304 = {1{`RANDOM}};
  _T_820_im = _RAND_1304[31:0];
  _RAND_1305 = {1{`RANDOM}};
  _T_821_re = _RAND_1305[31:0];
  _RAND_1306 = {1{`RANDOM}};
  _T_821_im = _RAND_1306[31:0];
  _RAND_1307 = {1{`RANDOM}};
  _T_822_re = _RAND_1307[31:0];
  _RAND_1308 = {1{`RANDOM}};
  _T_822_im = _RAND_1308[31:0];
  _RAND_1309 = {1{`RANDOM}};
  _T_823_re = _RAND_1309[31:0];
  _RAND_1310 = {1{`RANDOM}};
  _T_823_im = _RAND_1310[31:0];
  _RAND_1311 = {1{`RANDOM}};
  _T_824_re = _RAND_1311[31:0];
  _RAND_1312 = {1{`RANDOM}};
  _T_824_im = _RAND_1312[31:0];
  _RAND_1313 = {1{`RANDOM}};
  _T_825_re = _RAND_1313[31:0];
  _RAND_1314 = {1{`RANDOM}};
  _T_825_im = _RAND_1314[31:0];
  _RAND_1315 = {1{`RANDOM}};
  _T_826_re = _RAND_1315[31:0];
  _RAND_1316 = {1{`RANDOM}};
  _T_826_im = _RAND_1316[31:0];
  _RAND_1317 = {1{`RANDOM}};
  _T_827_re = _RAND_1317[31:0];
  _RAND_1318 = {1{`RANDOM}};
  _T_827_im = _RAND_1318[31:0];
  _RAND_1319 = {1{`RANDOM}};
  _T_828_re = _RAND_1319[31:0];
  _RAND_1320 = {1{`RANDOM}};
  _T_828_im = _RAND_1320[31:0];
  _RAND_1321 = {1{`RANDOM}};
  _T_829_re = _RAND_1321[31:0];
  _RAND_1322 = {1{`RANDOM}};
  _T_829_im = _RAND_1322[31:0];
  _RAND_1323 = {1{`RANDOM}};
  _T_830_re = _RAND_1323[31:0];
  _RAND_1324 = {1{`RANDOM}};
  _T_830_im = _RAND_1324[31:0];
  _RAND_1325 = {1{`RANDOM}};
  _T_831_re = _RAND_1325[31:0];
  _RAND_1326 = {1{`RANDOM}};
  _T_831_im = _RAND_1326[31:0];
  _RAND_1327 = {1{`RANDOM}};
  _T_832_re = _RAND_1327[31:0];
  _RAND_1328 = {1{`RANDOM}};
  _T_832_im = _RAND_1328[31:0];
  _RAND_1329 = {1{`RANDOM}};
  _T_833_re = _RAND_1329[31:0];
  _RAND_1330 = {1{`RANDOM}};
  _T_833_im = _RAND_1330[31:0];
  _RAND_1331 = {1{`RANDOM}};
  _T_834_re = _RAND_1331[31:0];
  _RAND_1332 = {1{`RANDOM}};
  _T_834_im = _RAND_1332[31:0];
  _RAND_1333 = {1{`RANDOM}};
  _T_835_re = _RAND_1333[31:0];
  _RAND_1334 = {1{`RANDOM}};
  _T_835_im = _RAND_1334[31:0];
  _RAND_1335 = {1{`RANDOM}};
  _T_836_re = _RAND_1335[31:0];
  _RAND_1336 = {1{`RANDOM}};
  _T_836_im = _RAND_1336[31:0];
  _RAND_1337 = {1{`RANDOM}};
  _T_837_re = _RAND_1337[31:0];
  _RAND_1338 = {1{`RANDOM}};
  _T_837_im = _RAND_1338[31:0];
  _RAND_1339 = {1{`RANDOM}};
  _T_838_re = _RAND_1339[31:0];
  _RAND_1340 = {1{`RANDOM}};
  _T_838_im = _RAND_1340[31:0];
  _RAND_1341 = {1{`RANDOM}};
  _T_839_re = _RAND_1341[31:0];
  _RAND_1342 = {1{`RANDOM}};
  _T_839_im = _RAND_1342[31:0];
  _RAND_1343 = {1{`RANDOM}};
  _T_840_re = _RAND_1343[31:0];
  _RAND_1344 = {1{`RANDOM}};
  _T_840_im = _RAND_1344[31:0];
  _RAND_1345 = {1{`RANDOM}};
  _T_849_re = _RAND_1345[31:0];
  _RAND_1346 = {1{`RANDOM}};
  _T_849_im = _RAND_1346[31:0];
  _RAND_1347 = {1{`RANDOM}};
  _T_850_re = _RAND_1347[31:0];
  _RAND_1348 = {1{`RANDOM}};
  _T_850_im = _RAND_1348[31:0];
  _RAND_1349 = {1{`RANDOM}};
  _T_851_re = _RAND_1349[31:0];
  _RAND_1350 = {1{`RANDOM}};
  _T_851_im = _RAND_1350[31:0];
  _RAND_1351 = {1{`RANDOM}};
  _T_852_re = _RAND_1351[31:0];
  _RAND_1352 = {1{`RANDOM}};
  _T_852_im = _RAND_1352[31:0];
  _RAND_1353 = {1{`RANDOM}};
  _T_853_re = _RAND_1353[31:0];
  _RAND_1354 = {1{`RANDOM}};
  _T_853_im = _RAND_1354[31:0];
  _RAND_1355 = {1{`RANDOM}};
  _T_854_re = _RAND_1355[31:0];
  _RAND_1356 = {1{`RANDOM}};
  _T_854_im = _RAND_1356[31:0];
  _RAND_1357 = {1{`RANDOM}};
  _T_855_re = _RAND_1357[31:0];
  _RAND_1358 = {1{`RANDOM}};
  _T_855_im = _RAND_1358[31:0];
  _RAND_1359 = {1{`RANDOM}};
  _T_856_re = _RAND_1359[31:0];
  _RAND_1360 = {1{`RANDOM}};
  _T_856_im = _RAND_1360[31:0];
  _RAND_1361 = {1{`RANDOM}};
  _T_857_re = _RAND_1361[31:0];
  _RAND_1362 = {1{`RANDOM}};
  _T_857_im = _RAND_1362[31:0];
  _RAND_1363 = {1{`RANDOM}};
  _T_858_re = _RAND_1363[31:0];
  _RAND_1364 = {1{`RANDOM}};
  _T_858_im = _RAND_1364[31:0];
  _RAND_1365 = {1{`RANDOM}};
  _T_859_re = _RAND_1365[31:0];
  _RAND_1366 = {1{`RANDOM}};
  _T_859_im = _RAND_1366[31:0];
  _RAND_1367 = {1{`RANDOM}};
  _T_860_re = _RAND_1367[31:0];
  _RAND_1368 = {1{`RANDOM}};
  _T_860_im = _RAND_1368[31:0];
  _RAND_1369 = {1{`RANDOM}};
  _T_861_re = _RAND_1369[31:0];
  _RAND_1370 = {1{`RANDOM}};
  _T_861_im = _RAND_1370[31:0];
  _RAND_1371 = {1{`RANDOM}};
  _T_862_re = _RAND_1371[31:0];
  _RAND_1372 = {1{`RANDOM}};
  _T_862_im = _RAND_1372[31:0];
  _RAND_1373 = {1{`RANDOM}};
  _T_863_re = _RAND_1373[31:0];
  _RAND_1374 = {1{`RANDOM}};
  _T_863_im = _RAND_1374[31:0];
  _RAND_1375 = {1{`RANDOM}};
  _T_864_re = _RAND_1375[31:0];
  _RAND_1376 = {1{`RANDOM}};
  _T_864_im = _RAND_1376[31:0];
  _RAND_1377 = {1{`RANDOM}};
  _T_865_re = _RAND_1377[31:0];
  _RAND_1378 = {1{`RANDOM}};
  _T_865_im = _RAND_1378[31:0];
  _RAND_1379 = {1{`RANDOM}};
  _T_866_re = _RAND_1379[31:0];
  _RAND_1380 = {1{`RANDOM}};
  _T_866_im = _RAND_1380[31:0];
  _RAND_1381 = {1{`RANDOM}};
  _T_867_re = _RAND_1381[31:0];
  _RAND_1382 = {1{`RANDOM}};
  _T_867_im = _RAND_1382[31:0];
  _RAND_1383 = {1{`RANDOM}};
  _T_868_re = _RAND_1383[31:0];
  _RAND_1384 = {1{`RANDOM}};
  _T_868_im = _RAND_1384[31:0];
  _RAND_1385 = {1{`RANDOM}};
  _T_869_re = _RAND_1385[31:0];
  _RAND_1386 = {1{`RANDOM}};
  _T_869_im = _RAND_1386[31:0];
  _RAND_1387 = {1{`RANDOM}};
  _T_870_re = _RAND_1387[31:0];
  _RAND_1388 = {1{`RANDOM}};
  _T_870_im = _RAND_1388[31:0];
  _RAND_1389 = {1{`RANDOM}};
  _T_871_re = _RAND_1389[31:0];
  _RAND_1390 = {1{`RANDOM}};
  _T_871_im = _RAND_1390[31:0];
  _RAND_1391 = {1{`RANDOM}};
  _T_872_re = _RAND_1391[31:0];
  _RAND_1392 = {1{`RANDOM}};
  _T_872_im = _RAND_1392[31:0];
  _RAND_1393 = {1{`RANDOM}};
  _T_873_re = _RAND_1393[31:0];
  _RAND_1394 = {1{`RANDOM}};
  _T_873_im = _RAND_1394[31:0];
  _RAND_1395 = {1{`RANDOM}};
  _T_874_re = _RAND_1395[31:0];
  _RAND_1396 = {1{`RANDOM}};
  _T_874_im = _RAND_1396[31:0];
  _RAND_1397 = {1{`RANDOM}};
  _T_875_re = _RAND_1397[31:0];
  _RAND_1398 = {1{`RANDOM}};
  _T_875_im = _RAND_1398[31:0];
  _RAND_1399 = {1{`RANDOM}};
  _T_876_re = _RAND_1399[31:0];
  _RAND_1400 = {1{`RANDOM}};
  _T_876_im = _RAND_1400[31:0];
  _RAND_1401 = {1{`RANDOM}};
  _T_877_re = _RAND_1401[31:0];
  _RAND_1402 = {1{`RANDOM}};
  _T_877_im = _RAND_1402[31:0];
  _RAND_1403 = {1{`RANDOM}};
  _T_878_re = _RAND_1403[31:0];
  _RAND_1404 = {1{`RANDOM}};
  _T_878_im = _RAND_1404[31:0];
  _RAND_1405 = {1{`RANDOM}};
  _T_879_re = _RAND_1405[31:0];
  _RAND_1406 = {1{`RANDOM}};
  _T_879_im = _RAND_1406[31:0];
  _RAND_1407 = {1{`RANDOM}};
  _T_880_re = _RAND_1407[31:0];
  _RAND_1408 = {1{`RANDOM}};
  _T_880_im = _RAND_1408[31:0];
  _RAND_1409 = {1{`RANDOM}};
  _T_882_re = _RAND_1409[31:0];
  _RAND_1410 = {1{`RANDOM}};
  _T_882_im = _RAND_1410[31:0];
  _RAND_1411 = {1{`RANDOM}};
  _T_883_re = _RAND_1411[31:0];
  _RAND_1412 = {1{`RANDOM}};
  _T_883_im = _RAND_1412[31:0];
  _RAND_1413 = {1{`RANDOM}};
  _T_884_re = _RAND_1413[31:0];
  _RAND_1414 = {1{`RANDOM}};
  _T_884_im = _RAND_1414[31:0];
  _RAND_1415 = {1{`RANDOM}};
  _T_885_re = _RAND_1415[31:0];
  _RAND_1416 = {1{`RANDOM}};
  _T_885_im = _RAND_1416[31:0];
  _RAND_1417 = {1{`RANDOM}};
  _T_886_re = _RAND_1417[31:0];
  _RAND_1418 = {1{`RANDOM}};
  _T_886_im = _RAND_1418[31:0];
  _RAND_1419 = {1{`RANDOM}};
  _T_887_re = _RAND_1419[31:0];
  _RAND_1420 = {1{`RANDOM}};
  _T_887_im = _RAND_1420[31:0];
  _RAND_1421 = {1{`RANDOM}};
  _T_888_re = _RAND_1421[31:0];
  _RAND_1422 = {1{`RANDOM}};
  _T_888_im = _RAND_1422[31:0];
  _RAND_1423 = {1{`RANDOM}};
  _T_889_re = _RAND_1423[31:0];
  _RAND_1424 = {1{`RANDOM}};
  _T_889_im = _RAND_1424[31:0];
  _RAND_1425 = {1{`RANDOM}};
  _T_890_re = _RAND_1425[31:0];
  _RAND_1426 = {1{`RANDOM}};
  _T_890_im = _RAND_1426[31:0];
  _RAND_1427 = {1{`RANDOM}};
  _T_891_re = _RAND_1427[31:0];
  _RAND_1428 = {1{`RANDOM}};
  _T_891_im = _RAND_1428[31:0];
  _RAND_1429 = {1{`RANDOM}};
  _T_892_re = _RAND_1429[31:0];
  _RAND_1430 = {1{`RANDOM}};
  _T_892_im = _RAND_1430[31:0];
  _RAND_1431 = {1{`RANDOM}};
  _T_893_re = _RAND_1431[31:0];
  _RAND_1432 = {1{`RANDOM}};
  _T_893_im = _RAND_1432[31:0];
  _RAND_1433 = {1{`RANDOM}};
  _T_894_re = _RAND_1433[31:0];
  _RAND_1434 = {1{`RANDOM}};
  _T_894_im = _RAND_1434[31:0];
  _RAND_1435 = {1{`RANDOM}};
  _T_895_re = _RAND_1435[31:0];
  _RAND_1436 = {1{`RANDOM}};
  _T_895_im = _RAND_1436[31:0];
  _RAND_1437 = {1{`RANDOM}};
  _T_896_re = _RAND_1437[31:0];
  _RAND_1438 = {1{`RANDOM}};
  _T_896_im = _RAND_1438[31:0];
  _RAND_1439 = {1{`RANDOM}};
  _T_897_re = _RAND_1439[31:0];
  _RAND_1440 = {1{`RANDOM}};
  _T_897_im = _RAND_1440[31:0];
  _RAND_1441 = {1{`RANDOM}};
  _T_906_re = _RAND_1441[31:0];
  _RAND_1442 = {1{`RANDOM}};
  _T_906_im = _RAND_1442[31:0];
  _RAND_1443 = {1{`RANDOM}};
  _T_907_re = _RAND_1443[31:0];
  _RAND_1444 = {1{`RANDOM}};
  _T_907_im = _RAND_1444[31:0];
  _RAND_1445 = {1{`RANDOM}};
  _T_908_re = _RAND_1445[31:0];
  _RAND_1446 = {1{`RANDOM}};
  _T_908_im = _RAND_1446[31:0];
  _RAND_1447 = {1{`RANDOM}};
  _T_909_re = _RAND_1447[31:0];
  _RAND_1448 = {1{`RANDOM}};
  _T_909_im = _RAND_1448[31:0];
  _RAND_1449 = {1{`RANDOM}};
  _T_910_re = _RAND_1449[31:0];
  _RAND_1450 = {1{`RANDOM}};
  _T_910_im = _RAND_1450[31:0];
  _RAND_1451 = {1{`RANDOM}};
  _T_911_re = _RAND_1451[31:0];
  _RAND_1452 = {1{`RANDOM}};
  _T_911_im = _RAND_1452[31:0];
  _RAND_1453 = {1{`RANDOM}};
  _T_912_re = _RAND_1453[31:0];
  _RAND_1454 = {1{`RANDOM}};
  _T_912_im = _RAND_1454[31:0];
  _RAND_1455 = {1{`RANDOM}};
  _T_913_re = _RAND_1455[31:0];
  _RAND_1456 = {1{`RANDOM}};
  _T_913_im = _RAND_1456[31:0];
  _RAND_1457 = {1{`RANDOM}};
  _T_914_re = _RAND_1457[31:0];
  _RAND_1458 = {1{`RANDOM}};
  _T_914_im = _RAND_1458[31:0];
  _RAND_1459 = {1{`RANDOM}};
  _T_915_re = _RAND_1459[31:0];
  _RAND_1460 = {1{`RANDOM}};
  _T_915_im = _RAND_1460[31:0];
  _RAND_1461 = {1{`RANDOM}};
  _T_916_re = _RAND_1461[31:0];
  _RAND_1462 = {1{`RANDOM}};
  _T_916_im = _RAND_1462[31:0];
  _RAND_1463 = {1{`RANDOM}};
  _T_917_re = _RAND_1463[31:0];
  _RAND_1464 = {1{`RANDOM}};
  _T_917_im = _RAND_1464[31:0];
  _RAND_1465 = {1{`RANDOM}};
  _T_918_re = _RAND_1465[31:0];
  _RAND_1466 = {1{`RANDOM}};
  _T_918_im = _RAND_1466[31:0];
  _RAND_1467 = {1{`RANDOM}};
  _T_919_re = _RAND_1467[31:0];
  _RAND_1468 = {1{`RANDOM}};
  _T_919_im = _RAND_1468[31:0];
  _RAND_1469 = {1{`RANDOM}};
  _T_920_re = _RAND_1469[31:0];
  _RAND_1470 = {1{`RANDOM}};
  _T_920_im = _RAND_1470[31:0];
  _RAND_1471 = {1{`RANDOM}};
  _T_921_re = _RAND_1471[31:0];
  _RAND_1472 = {1{`RANDOM}};
  _T_921_im = _RAND_1472[31:0];
  _RAND_1473 = {1{`RANDOM}};
  _T_923_re = _RAND_1473[31:0];
  _RAND_1474 = {1{`RANDOM}};
  _T_923_im = _RAND_1474[31:0];
  _RAND_1475 = {1{`RANDOM}};
  _T_924_re = _RAND_1475[31:0];
  _RAND_1476 = {1{`RANDOM}};
  _T_924_im = _RAND_1476[31:0];
  _RAND_1477 = {1{`RANDOM}};
  _T_925_re = _RAND_1477[31:0];
  _RAND_1478 = {1{`RANDOM}};
  _T_925_im = _RAND_1478[31:0];
  _RAND_1479 = {1{`RANDOM}};
  _T_926_re = _RAND_1479[31:0];
  _RAND_1480 = {1{`RANDOM}};
  _T_926_im = _RAND_1480[31:0];
  _RAND_1481 = {1{`RANDOM}};
  _T_927_re = _RAND_1481[31:0];
  _RAND_1482 = {1{`RANDOM}};
  _T_927_im = _RAND_1482[31:0];
  _RAND_1483 = {1{`RANDOM}};
  _T_928_re = _RAND_1483[31:0];
  _RAND_1484 = {1{`RANDOM}};
  _T_928_im = _RAND_1484[31:0];
  _RAND_1485 = {1{`RANDOM}};
  _T_929_re = _RAND_1485[31:0];
  _RAND_1486 = {1{`RANDOM}};
  _T_929_im = _RAND_1486[31:0];
  _RAND_1487 = {1{`RANDOM}};
  _T_930_re = _RAND_1487[31:0];
  _RAND_1488 = {1{`RANDOM}};
  _T_930_im = _RAND_1488[31:0];
  _RAND_1489 = {1{`RANDOM}};
  _T_939_re = _RAND_1489[31:0];
  _RAND_1490 = {1{`RANDOM}};
  _T_939_im = _RAND_1490[31:0];
  _RAND_1491 = {1{`RANDOM}};
  _T_940_re = _RAND_1491[31:0];
  _RAND_1492 = {1{`RANDOM}};
  _T_940_im = _RAND_1492[31:0];
  _RAND_1493 = {1{`RANDOM}};
  _T_941_re = _RAND_1493[31:0];
  _RAND_1494 = {1{`RANDOM}};
  _T_941_im = _RAND_1494[31:0];
  _RAND_1495 = {1{`RANDOM}};
  _T_942_re = _RAND_1495[31:0];
  _RAND_1496 = {1{`RANDOM}};
  _T_942_im = _RAND_1496[31:0];
  _RAND_1497 = {1{`RANDOM}};
  _T_943_re = _RAND_1497[31:0];
  _RAND_1498 = {1{`RANDOM}};
  _T_943_im = _RAND_1498[31:0];
  _RAND_1499 = {1{`RANDOM}};
  _T_944_re = _RAND_1499[31:0];
  _RAND_1500 = {1{`RANDOM}};
  _T_944_im = _RAND_1500[31:0];
  _RAND_1501 = {1{`RANDOM}};
  _T_945_re = _RAND_1501[31:0];
  _RAND_1502 = {1{`RANDOM}};
  _T_945_im = _RAND_1502[31:0];
  _RAND_1503 = {1{`RANDOM}};
  _T_946_re = _RAND_1503[31:0];
  _RAND_1504 = {1{`RANDOM}};
  _T_946_im = _RAND_1504[31:0];
  _RAND_1505 = {1{`RANDOM}};
  _T_948_re = _RAND_1505[31:0];
  _RAND_1506 = {1{`RANDOM}};
  _T_948_im = _RAND_1506[31:0];
  _RAND_1507 = {1{`RANDOM}};
  _T_949_re = _RAND_1507[31:0];
  _RAND_1508 = {1{`RANDOM}};
  _T_949_im = _RAND_1508[31:0];
  _RAND_1509 = {1{`RANDOM}};
  _T_950_re = _RAND_1509[31:0];
  _RAND_1510 = {1{`RANDOM}};
  _T_950_im = _RAND_1510[31:0];
  _RAND_1511 = {1{`RANDOM}};
  _T_951_re = _RAND_1511[31:0];
  _RAND_1512 = {1{`RANDOM}};
  _T_951_im = _RAND_1512[31:0];
  _RAND_1513 = {1{`RANDOM}};
  _T_960_re = _RAND_1513[31:0];
  _RAND_1514 = {1{`RANDOM}};
  _T_960_im = _RAND_1514[31:0];
  _RAND_1515 = {1{`RANDOM}};
  _T_961_re = _RAND_1515[31:0];
  _RAND_1516 = {1{`RANDOM}};
  _T_961_im = _RAND_1516[31:0];
  _RAND_1517 = {1{`RANDOM}};
  _T_962_re = _RAND_1517[31:0];
  _RAND_1518 = {1{`RANDOM}};
  _T_962_im = _RAND_1518[31:0];
  _RAND_1519 = {1{`RANDOM}};
  _T_963_re = _RAND_1519[31:0];
  _RAND_1520 = {1{`RANDOM}};
  _T_963_im = _RAND_1520[31:0];
  _RAND_1521 = {1{`RANDOM}};
  _T_965_re = _RAND_1521[31:0];
  _RAND_1522 = {1{`RANDOM}};
  _T_965_im = _RAND_1522[31:0];
  _RAND_1523 = {1{`RANDOM}};
  _T_966_re = _RAND_1523[31:0];
  _RAND_1524 = {1{`RANDOM}};
  _T_966_im = _RAND_1524[31:0];
  _RAND_1525 = {1{`RANDOM}};
  _T_975_re = _RAND_1525[31:0];
  _RAND_1526 = {1{`RANDOM}};
  _T_975_im = _RAND_1526[31:0];
  _RAND_1527 = {1{`RANDOM}};
  _T_976_re = _RAND_1527[31:0];
  _RAND_1528 = {1{`RANDOM}};
  _T_976_im = _RAND_1528[31:0];
  _RAND_1529 = {1{`RANDOM}};
  _T_978_re = _RAND_1529[31:0];
  _RAND_1530 = {1{`RANDOM}};
  _T_978_im = _RAND_1530[31:0];
  _RAND_1531 = {1{`RANDOM}};
  out1D1_re = _RAND_1531[31:0];
  _RAND_1532 = {1{`RANDOM}};
  out1D1_im = _RAND_1532[31:0];
  _RAND_1533 = {1{`RANDOM}};
  _T_985_re = _RAND_1533[31:0];
  _RAND_1534 = {1{`RANDOM}};
  _T_985_im = _RAND_1534[31:0];
  _RAND_1535 = {1{`RANDOM}};
  _T_986_re = _RAND_1535[31:0];
  _RAND_1536 = {1{`RANDOM}};
  _T_986_im = _RAND_1536[31:0];
  _RAND_1537 = {1{`RANDOM}};
  _T_987 = _RAND_1537[0:0];
  _RAND_1538 = {1{`RANDOM}};
  _T_988 = _RAND_1538[0:0];
  _RAND_1539 = {1{`RANDOM}};
  _T_989 = _RAND_1539[0:0];
  _RAND_1540 = {1{`RANDOM}};
  _T_990 = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  _T_991 = _RAND_1541[0:0];
  _RAND_1542 = {1{`RANDOM}};
  _T_992 = _RAND_1542[0:0];
  _RAND_1543 = {1{`RANDOM}};
  _T_993 = _RAND_1543[0:0];
  _RAND_1544 = {1{`RANDOM}};
  _T_994 = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  _T_995 = _RAND_1545[0:0];
  _RAND_1546 = {1{`RANDOM}};
  _T_996 = _RAND_1546[0:0];
  _RAND_1547 = {1{`RANDOM}};
  _T_997 = _RAND_1547[0:0];
  _RAND_1548 = {1{`RANDOM}};
  _T_998 = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  _T_999 = _RAND_1549[0:0];
  _RAND_1550 = {1{`RANDOM}};
  _T_1000 = _RAND_1550[0:0];
  _RAND_1551 = {1{`RANDOM}};
  _T_1001 = _RAND_1551[0:0];
  _RAND_1552 = {1{`RANDOM}};
  _T_1002 = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  _T_1003 = _RAND_1553[0:0];
  _RAND_1554 = {1{`RANDOM}};
  _T_1004 = _RAND_1554[0:0];
  _RAND_1555 = {1{`RANDOM}};
  _T_1005 = _RAND_1555[0:0];
  _RAND_1556 = {1{`RANDOM}};
  _T_1006 = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  _T_1007 = _RAND_1557[0:0];
  _RAND_1558 = {1{`RANDOM}};
  _T_1008 = _RAND_1558[0:0];
  _RAND_1559 = {1{`RANDOM}};
  _T_1009 = _RAND_1559[0:0];
  _RAND_1560 = {1{`RANDOM}};
  _T_1010 = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  _T_1011 = _RAND_1561[0:0];
  _RAND_1562 = {1{`RANDOM}};
  _T_1012 = _RAND_1562[0:0];
  _RAND_1563 = {1{`RANDOM}};
  _T_1013 = _RAND_1563[0:0];
  _RAND_1564 = {1{`RANDOM}};
  _T_1014 = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  _T_1015 = _RAND_1565[0:0];
  _RAND_1566 = {1{`RANDOM}};
  _T_1016 = _RAND_1566[0:0];
  _RAND_1567 = {1{`RANDOM}};
  _T_1017 = _RAND_1567[0:0];
  _RAND_1568 = {1{`RANDOM}};
  _T_1018 = _RAND_1568[0:0];
  _RAND_1569 = {1{`RANDOM}};
  _T_1019 = _RAND_1569[0:0];
  _RAND_1570 = {1{`RANDOM}};
  _T_1020 = _RAND_1570[0:0];
  _RAND_1571 = {1{`RANDOM}};
  _T_1021 = _RAND_1571[0:0];
  _RAND_1572 = {1{`RANDOM}};
  _T_1022 = _RAND_1572[0:0];
  _RAND_1573 = {1{`RANDOM}};
  _T_1023 = _RAND_1573[0:0];
  _RAND_1574 = {1{`RANDOM}};
  _T_1024 = _RAND_1574[0:0];
  _RAND_1575 = {1{`RANDOM}};
  _T_1025 = _RAND_1575[0:0];
  _RAND_1576 = {1{`RANDOM}};
  _T_1026 = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  _T_1027 = _RAND_1577[0:0];
  _RAND_1578 = {1{`RANDOM}};
  _T_1028 = _RAND_1578[0:0];
  _RAND_1579 = {1{`RANDOM}};
  _T_1029 = _RAND_1579[0:0];
  _RAND_1580 = {1{`RANDOM}};
  _T_1030 = _RAND_1580[0:0];
  _RAND_1581 = {1{`RANDOM}};
  _T_1031 = _RAND_1581[0:0];
  _RAND_1582 = {1{`RANDOM}};
  _T_1032 = _RAND_1582[0:0];
  _RAND_1583 = {1{`RANDOM}};
  _T_1033 = _RAND_1583[0:0];
  _RAND_1584 = {1{`RANDOM}};
  _T_1034 = _RAND_1584[0:0];
  _RAND_1585 = {1{`RANDOM}};
  _T_1035 = _RAND_1585[0:0];
  _RAND_1586 = {1{`RANDOM}};
  _T_1036 = _RAND_1586[0:0];
  _RAND_1587 = {1{`RANDOM}};
  _T_1037 = _RAND_1587[0:0];
  _RAND_1588 = {1{`RANDOM}};
  _T_1038 = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  _T_1039 = _RAND_1589[0:0];
  _RAND_1590 = {1{`RANDOM}};
  _T_1040 = _RAND_1590[0:0];
  _RAND_1591 = {1{`RANDOM}};
  _T_1041 = _RAND_1591[0:0];
  _RAND_1592 = {1{`RANDOM}};
  _T_1042 = _RAND_1592[0:0];
  _RAND_1593 = {1{`RANDOM}};
  _T_1043 = _RAND_1593[0:0];
  _RAND_1594 = {1{`RANDOM}};
  _T_1044 = _RAND_1594[0:0];
  _RAND_1595 = {1{`RANDOM}};
  _T_1045 = _RAND_1595[0:0];
  _RAND_1596 = {1{`RANDOM}};
  _T_1046 = _RAND_1596[0:0];
  _RAND_1597 = {1{`RANDOM}};
  _T_1047 = _RAND_1597[0:0];
  _RAND_1598 = {1{`RANDOM}};
  _T_1048 = _RAND_1598[0:0];
  _RAND_1599 = {1{`RANDOM}};
  _T_1049 = _RAND_1599[0:0];
  _RAND_1600 = {1{`RANDOM}};
  _T_1050 = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  _T_1051 = _RAND_1601[0:0];
  _RAND_1602 = {1{`RANDOM}};
  _T_1052 = _RAND_1602[0:0];
  _RAND_1603 = {1{`RANDOM}};
  _T_1053 = _RAND_1603[0:0];
  _RAND_1604 = {1{`RANDOM}};
  _T_1054 = _RAND_1604[0:0];
  _RAND_1605 = {1{`RANDOM}};
  _T_1055 = _RAND_1605[0:0];
  _RAND_1606 = {1{`RANDOM}};
  _T_1056 = _RAND_1606[0:0];
  _RAND_1607 = {1{`RANDOM}};
  _T_1057 = _RAND_1607[0:0];
  _RAND_1608 = {1{`RANDOM}};
  _T_1058 = _RAND_1608[0:0];
  _RAND_1609 = {1{`RANDOM}};
  _T_1059 = _RAND_1609[0:0];
  _RAND_1610 = {1{`RANDOM}};
  _T_1060 = _RAND_1610[0:0];
  _RAND_1611 = {1{`RANDOM}};
  _T_1061 = _RAND_1611[0:0];
  _RAND_1612 = {1{`RANDOM}};
  _T_1062 = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  _T_1063 = _RAND_1613[0:0];
  _RAND_1614 = {1{`RANDOM}};
  _T_1064 = _RAND_1614[0:0];
  _RAND_1615 = {1{`RANDOM}};
  _T_1065 = _RAND_1615[0:0];
  _RAND_1616 = {1{`RANDOM}};
  _T_1066 = _RAND_1616[0:0];
  _RAND_1617 = {1{`RANDOM}};
  _T_1067 = _RAND_1617[0:0];
  _RAND_1618 = {1{`RANDOM}};
  _T_1068 = _RAND_1618[0:0];
  _RAND_1619 = {1{`RANDOM}};
  _T_1069 = _RAND_1619[0:0];
  _RAND_1620 = {1{`RANDOM}};
  _T_1070 = _RAND_1620[0:0];
  _RAND_1621 = {1{`RANDOM}};
  _T_1071 = _RAND_1621[0:0];
  _RAND_1622 = {1{`RANDOM}};
  _T_1072 = _RAND_1622[0:0];
  _RAND_1623 = {1{`RANDOM}};
  _T_1073 = _RAND_1623[0:0];
  _RAND_1624 = {1{`RANDOM}};
  _T_1074 = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  _T_1075 = _RAND_1625[0:0];
  _RAND_1626 = {1{`RANDOM}};
  _T_1076 = _RAND_1626[0:0];
  _RAND_1627 = {1{`RANDOM}};
  _T_1077 = _RAND_1627[0:0];
  _RAND_1628 = {1{`RANDOM}};
  _T_1078 = _RAND_1628[0:0];
  _RAND_1629 = {1{`RANDOM}};
  _T_1079 = _RAND_1629[0:0];
  _RAND_1630 = {1{`RANDOM}};
  _T_1080 = _RAND_1630[0:0];
  _RAND_1631 = {1{`RANDOM}};
  _T_1081 = _RAND_1631[0:0];
  _RAND_1632 = {1{`RANDOM}};
  _T_1082 = _RAND_1632[0:0];
  _RAND_1633 = {1{`RANDOM}};
  _T_1083 = _RAND_1633[0:0];
  _RAND_1634 = {1{`RANDOM}};
  _T_1084 = _RAND_1634[0:0];
  _RAND_1635 = {1{`RANDOM}};
  _T_1085 = _RAND_1635[0:0];
  _RAND_1636 = {1{`RANDOM}};
  _T_1086 = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  _T_1087 = _RAND_1637[0:0];
  _RAND_1638 = {1{`RANDOM}};
  _T_1088 = _RAND_1638[0:0];
  _RAND_1639 = {1{`RANDOM}};
  _T_1089 = _RAND_1639[0:0];
  _RAND_1640 = {1{`RANDOM}};
  _T_1090 = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  _T_1091 = _RAND_1641[0:0];
  _RAND_1642 = {1{`RANDOM}};
  _T_1092 = _RAND_1642[0:0];
  _RAND_1643 = {1{`RANDOM}};
  _T_1093 = _RAND_1643[0:0];
  _RAND_1644 = {1{`RANDOM}};
  _T_1094 = _RAND_1644[0:0];
  _RAND_1645 = {1{`RANDOM}};
  _T_1095 = _RAND_1645[0:0];
  _RAND_1646 = {1{`RANDOM}};
  _T_1096 = _RAND_1646[0:0];
  _RAND_1647 = {1{`RANDOM}};
  _T_1097 = _RAND_1647[0:0];
  _RAND_1648 = {1{`RANDOM}};
  _T_1098 = _RAND_1648[0:0];
  _RAND_1649 = {1{`RANDOM}};
  _T_1099 = _RAND_1649[0:0];
  _RAND_1650 = {1{`RANDOM}};
  _T_1100 = _RAND_1650[0:0];
  _RAND_1651 = {1{`RANDOM}};
  _T_1101 = _RAND_1651[0:0];
  _RAND_1652 = {1{`RANDOM}};
  _T_1102 = _RAND_1652[0:0];
  _RAND_1653 = {1{`RANDOM}};
  _T_1103 = _RAND_1653[0:0];
  _RAND_1654 = {1{`RANDOM}};
  _T_1104 = _RAND_1654[0:0];
  _RAND_1655 = {1{`RANDOM}};
  _T_1105 = _RAND_1655[0:0];
  _RAND_1656 = {1{`RANDOM}};
  _T_1106 = _RAND_1656[0:0];
  _RAND_1657 = {1{`RANDOM}};
  _T_1107 = _RAND_1657[0:0];
  _RAND_1658 = {1{`RANDOM}};
  _T_1108 = _RAND_1658[0:0];
  _RAND_1659 = {1{`RANDOM}};
  _T_1109 = _RAND_1659[0:0];
  _RAND_1660 = {1{`RANDOM}};
  _T_1110 = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  _T_1111 = _RAND_1661[0:0];
  _RAND_1662 = {1{`RANDOM}};
  _T_1112 = _RAND_1662[0:0];
  _RAND_1663 = {1{`RANDOM}};
  _T_1113 = _RAND_1663[0:0];
  _RAND_1664 = {1{`RANDOM}};
  _T_1114 = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  _T_1115 = _RAND_1665[0:0];
  _RAND_1666 = {1{`RANDOM}};
  _T_1116 = _RAND_1666[0:0];
  _RAND_1667 = {1{`RANDOM}};
  _T_1117 = _RAND_1667[0:0];
  _RAND_1668 = {1{`RANDOM}};
  _T_1118 = _RAND_1668[0:0];
  _RAND_1669 = {1{`RANDOM}};
  _T_1119 = _RAND_1669[0:0];
  _RAND_1670 = {1{`RANDOM}};
  _T_1120 = _RAND_1670[0:0];
  _RAND_1671 = {1{`RANDOM}};
  _T_1121 = _RAND_1671[0:0];
  _RAND_1672 = {1{`RANDOM}};
  _T_1122 = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  _T_1123 = _RAND_1673[0:0];
  _RAND_1674 = {1{`RANDOM}};
  _T_1124 = _RAND_1674[0:0];
  _RAND_1675 = {1{`RANDOM}};
  _T_1125 = _RAND_1675[0:0];
  _RAND_1676 = {1{`RANDOM}};
  _T_1126 = _RAND_1676[0:0];
  _RAND_1677 = {1{`RANDOM}};
  _T_1127 = _RAND_1677[0:0];
  _RAND_1678 = {1{`RANDOM}};
  _T_1128 = _RAND_1678[0:0];
  _RAND_1679 = {1{`RANDOM}};
  _T_1129 = _RAND_1679[0:0];
  _RAND_1680 = {1{`RANDOM}};
  _T_1130 = _RAND_1680[0:0];
  _RAND_1681 = {1{`RANDOM}};
  _T_1131 = _RAND_1681[0:0];
  _RAND_1682 = {1{`RANDOM}};
  _T_1132 = _RAND_1682[0:0];
  _RAND_1683 = {1{`RANDOM}};
  _T_1133 = _RAND_1683[0:0];
  _RAND_1684 = {1{`RANDOM}};
  _T_1134 = _RAND_1684[0:0];
  _RAND_1685 = {1{`RANDOM}};
  _T_1135 = _RAND_1685[0:0];
  _RAND_1686 = {1{`RANDOM}};
  _T_1136 = _RAND_1686[0:0];
  _RAND_1687 = {1{`RANDOM}};
  _T_1137 = _RAND_1687[0:0];
  _RAND_1688 = {1{`RANDOM}};
  _T_1138 = _RAND_1688[0:0];
  _RAND_1689 = {1{`RANDOM}};
  _T_1139 = _RAND_1689[0:0];
  _RAND_1690 = {1{`RANDOM}};
  _T_1140 = _RAND_1690[0:0];
  _RAND_1691 = {1{`RANDOM}};
  _T_1141 = _RAND_1691[0:0];
  _RAND_1692 = {1{`RANDOM}};
  _T_1142 = _RAND_1692[0:0];
  _RAND_1693 = {1{`RANDOM}};
  _T_1143 = _RAND_1693[0:0];
  _RAND_1694 = {1{`RANDOM}};
  _T_1144 = _RAND_1694[0:0];
  _RAND_1695 = {1{`RANDOM}};
  _T_1145 = _RAND_1695[0:0];
  _RAND_1696 = {1{`RANDOM}};
  _T_1146 = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  _T_1147 = _RAND_1697[0:0];
  _RAND_1698 = {1{`RANDOM}};
  _T_1148 = _RAND_1698[0:0];
  _RAND_1699 = {1{`RANDOM}};
  _T_1149 = _RAND_1699[0:0];
  _RAND_1700 = {1{`RANDOM}};
  _T_1150 = _RAND_1700[0:0];
  _RAND_1701 = {1{`RANDOM}};
  _T_1151 = _RAND_1701[0:0];
  _RAND_1702 = {1{`RANDOM}};
  _T_1152 = _RAND_1702[0:0];
  _RAND_1703 = {1{`RANDOM}};
  _T_1153 = _RAND_1703[0:0];
  _RAND_1704 = {1{`RANDOM}};
  _T_1154 = _RAND_1704[0:0];
  _RAND_1705 = {1{`RANDOM}};
  _T_1155 = _RAND_1705[0:0];
  _RAND_1706 = {1{`RANDOM}};
  _T_1156 = _RAND_1706[0:0];
  _RAND_1707 = {1{`RANDOM}};
  _T_1157 = _RAND_1707[0:0];
  _RAND_1708 = {1{`RANDOM}};
  _T_1158 = _RAND_1708[0:0];
  _RAND_1709 = {1{`RANDOM}};
  _T_1159 = _RAND_1709[0:0];
  _RAND_1710 = {1{`RANDOM}};
  _T_1160 = _RAND_1710[0:0];
  _RAND_1711 = {1{`RANDOM}};
  _T_1161 = _RAND_1711[0:0];
  _RAND_1712 = {1{`RANDOM}};
  _T_1162 = _RAND_1712[0:0];
  _RAND_1713 = {1{`RANDOM}};
  _T_1163 = _RAND_1713[0:0];
  _RAND_1714 = {1{`RANDOM}};
  _T_1164 = _RAND_1714[0:0];
  _RAND_1715 = {1{`RANDOM}};
  _T_1165 = _RAND_1715[0:0];
  _RAND_1716 = {1{`RANDOM}};
  _T_1166 = _RAND_1716[0:0];
  _RAND_1717 = {1{`RANDOM}};
  _T_1167 = _RAND_1717[0:0];
  _RAND_1718 = {1{`RANDOM}};
  _T_1168 = _RAND_1718[0:0];
  _RAND_1719 = {1{`RANDOM}};
  _T_1169 = _RAND_1719[0:0];
  _RAND_1720 = {1{`RANDOM}};
  _T_1170 = _RAND_1720[0:0];
  _RAND_1721 = {1{`RANDOM}};
  _T_1171 = _RAND_1721[0:0];
  _RAND_1722 = {1{`RANDOM}};
  _T_1172 = _RAND_1722[0:0];
  _RAND_1723 = {1{`RANDOM}};
  _T_1173 = _RAND_1723[0:0];
  _RAND_1724 = {1{`RANDOM}};
  _T_1174 = _RAND_1724[0:0];
  _RAND_1725 = {1{`RANDOM}};
  _T_1175 = _RAND_1725[0:0];
  _RAND_1726 = {1{`RANDOM}};
  _T_1176 = _RAND_1726[0:0];
  _RAND_1727 = {1{`RANDOM}};
  _T_1177 = _RAND_1727[0:0];
  _RAND_1728 = {1{`RANDOM}};
  _T_1178 = _RAND_1728[0:0];
  _RAND_1729 = {1{`RANDOM}};
  _T_1179 = _RAND_1729[0:0];
  _RAND_1730 = {1{`RANDOM}};
  _T_1180 = _RAND_1730[0:0];
  _RAND_1731 = {1{`RANDOM}};
  _T_1181 = _RAND_1731[0:0];
  _RAND_1732 = {1{`RANDOM}};
  _T_1182 = _RAND_1732[0:0];
  _RAND_1733 = {1{`RANDOM}};
  _T_1183 = _RAND_1733[0:0];
  _RAND_1734 = {1{`RANDOM}};
  _T_1184 = _RAND_1734[0:0];
  _RAND_1735 = {1{`RANDOM}};
  _T_1185 = _RAND_1735[0:0];
  _RAND_1736 = {1{`RANDOM}};
  _T_1186 = _RAND_1736[0:0];
  _RAND_1737 = {1{`RANDOM}};
  _T_1187 = _RAND_1737[0:0];
  _RAND_1738 = {1{`RANDOM}};
  _T_1188 = _RAND_1738[0:0];
  _RAND_1739 = {1{`RANDOM}};
  _T_1189 = _RAND_1739[0:0];
  _RAND_1740 = {1{`RANDOM}};
  _T_1190 = _RAND_1740[0:0];
  _RAND_1741 = {1{`RANDOM}};
  _T_1191 = _RAND_1741[0:0];
  _RAND_1742 = {1{`RANDOM}};
  _T_1192 = _RAND_1742[0:0];
  _RAND_1743 = {1{`RANDOM}};
  _T_1193 = _RAND_1743[0:0];
  _RAND_1744 = {1{`RANDOM}};
  _T_1194 = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  _T_1195 = _RAND_1745[0:0];
  _RAND_1746 = {1{`RANDOM}};
  _T_1196 = _RAND_1746[0:0];
  _RAND_1747 = {1{`RANDOM}};
  _T_1197 = _RAND_1747[0:0];
  _RAND_1748 = {1{`RANDOM}};
  _T_1198 = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  _T_1199 = _RAND_1749[0:0];
  _RAND_1750 = {1{`RANDOM}};
  _T_1200 = _RAND_1750[0:0];
  _RAND_1751 = {1{`RANDOM}};
  _T_1201 = _RAND_1751[0:0];
  _RAND_1752 = {1{`RANDOM}};
  _T_1202 = _RAND_1752[0:0];
  _RAND_1753 = {1{`RANDOM}};
  _T_1203 = _RAND_1753[0:0];
  _RAND_1754 = {1{`RANDOM}};
  _T_1204 = _RAND_1754[0:0];
  _RAND_1755 = {1{`RANDOM}};
  _T_1205 = _RAND_1755[0:0];
  _RAND_1756 = {1{`RANDOM}};
  _T_1206 = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  _T_1207 = _RAND_1757[0:0];
  _RAND_1758 = {1{`RANDOM}};
  _T_1208 = _RAND_1758[0:0];
  _RAND_1759 = {1{`RANDOM}};
  _T_1209 = _RAND_1759[0:0];
  _RAND_1760 = {1{`RANDOM}};
  _T_1210 = _RAND_1760[0:0];
  _RAND_1761 = {1{`RANDOM}};
  _T_1211 = _RAND_1761[0:0];
  _RAND_1762 = {1{`RANDOM}};
  _T_1212 = _RAND_1762[0:0];
  _RAND_1763 = {1{`RANDOM}};
  _T_1213 = _RAND_1763[0:0];
  _RAND_1764 = {1{`RANDOM}};
  _T_1214 = _RAND_1764[0:0];
  _RAND_1765 = {1{`RANDOM}};
  _T_1215 = _RAND_1765[0:0];
  _RAND_1766 = {1{`RANDOM}};
  _T_1216 = _RAND_1766[0:0];
  _RAND_1767 = {1{`RANDOM}};
  _T_1217 = _RAND_1767[0:0];
  _RAND_1768 = {1{`RANDOM}};
  _T_1218 = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  _T_1219 = _RAND_1769[0:0];
  _RAND_1770 = {1{`RANDOM}};
  _T_1220 = _RAND_1770[0:0];
  _RAND_1771 = {1{`RANDOM}};
  _T_1221 = _RAND_1771[0:0];
  _RAND_1772 = {1{`RANDOM}};
  _T_1222 = _RAND_1772[0:0];
  _RAND_1773 = {1{`RANDOM}};
  _T_1223 = _RAND_1773[0:0];
  _RAND_1774 = {1{`RANDOM}};
  _T_1224 = _RAND_1774[0:0];
  _RAND_1775 = {1{`RANDOM}};
  _T_1225 = _RAND_1775[0:0];
  _RAND_1776 = {1{`RANDOM}};
  _T_1226 = _RAND_1776[0:0];
  _RAND_1777 = {1{`RANDOM}};
  _T_1227 = _RAND_1777[0:0];
  _RAND_1778 = {1{`RANDOM}};
  _T_1228 = _RAND_1778[0:0];
  _RAND_1779 = {1{`RANDOM}};
  _T_1229 = _RAND_1779[0:0];
  _RAND_1780 = {1{`RANDOM}};
  _T_1230 = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  _T_1231 = _RAND_1781[0:0];
  _RAND_1782 = {1{`RANDOM}};
  _T_1232 = _RAND_1782[0:0];
  _RAND_1783 = {1{`RANDOM}};
  _T_1233 = _RAND_1783[0:0];
  _RAND_1784 = {1{`RANDOM}};
  _T_1234 = _RAND_1784[0:0];
  _RAND_1785 = {1{`RANDOM}};
  _T_1235 = _RAND_1785[0:0];
  _RAND_1786 = {1{`RANDOM}};
  _T_1236 = _RAND_1786[0:0];
  _RAND_1787 = {1{`RANDOM}};
  _T_1237 = _RAND_1787[0:0];
  _RAND_1788 = {1{`RANDOM}};
  _T_1238 = _RAND_1788[0:0];
  _RAND_1789 = {1{`RANDOM}};
  _T_1239 = _RAND_1789[0:0];
  _RAND_1790 = {1{`RANDOM}};
  _T_1240 = _RAND_1790[0:0];
  _RAND_1791 = {1{`RANDOM}};
  _T_1241 = _RAND_1791[0:0];
  _RAND_1792 = {1{`RANDOM}};
  _T_1242 = _RAND_1792[0:0];
  _RAND_1793 = {1{`RANDOM}};
  _T_1243 = _RAND_1793[0:0];
  _RAND_1794 = {1{`RANDOM}};
  _T_1244 = _RAND_1794[0:0];
  _RAND_1795 = {1{`RANDOM}};
  _T_1245 = _RAND_1795[0:0];
  _RAND_1796 = {1{`RANDOM}};
  _T_1246 = _RAND_1796[0:0];
  _RAND_1797 = {1{`RANDOM}};
  _T_1247 = _RAND_1797[0:0];
  _RAND_1798 = {1{`RANDOM}};
  _T_1248 = _RAND_1798[0:0];
  _RAND_1799 = {1{`RANDOM}};
  _T_1249 = _RAND_1799[0:0];
  _RAND_1800 = {1{`RANDOM}};
  _T_1250 = _RAND_1800[0:0];
  _RAND_1801 = {1{`RANDOM}};
  _T_1251 = _RAND_1801[0:0];
  _RAND_1802 = {1{`RANDOM}};
  _T_1252 = _RAND_1802[0:0];
  _RAND_1803 = {1{`RANDOM}};
  _T_1253 = _RAND_1803[0:0];
  _RAND_1804 = {1{`RANDOM}};
  _T_1254 = _RAND_1804[0:0];
  _RAND_1805 = {1{`RANDOM}};
  _T_1255 = _RAND_1805[0:0];
  _RAND_1806 = {1{`RANDOM}};
  _T_1256 = _RAND_1806[0:0];
  _RAND_1807 = {1{`RANDOM}};
  _T_1257 = _RAND_1807[0:0];
  _RAND_1808 = {1{`RANDOM}};
  _T_1258 = _RAND_1808[0:0];
  _RAND_1809 = {1{`RANDOM}};
  _T_1259 = _RAND_1809[0:0];
  _RAND_1810 = {1{`RANDOM}};
  _T_1260 = _RAND_1810[0:0];
  _RAND_1811 = {1{`RANDOM}};
  _T_1261 = _RAND_1811[0:0];
  _RAND_1812 = {1{`RANDOM}};
  _T_1262 = _RAND_1812[0:0];
  _RAND_1813 = {1{`RANDOM}};
  _T_1263 = _RAND_1813[0:0];
  _RAND_1814 = {1{`RANDOM}};
  _T_1264 = _RAND_1814[0:0];
  _RAND_1815 = {1{`RANDOM}};
  _T_1265 = _RAND_1815[0:0];
  _RAND_1816 = {1{`RANDOM}};
  _T_1266 = _RAND_1816[0:0];
  _RAND_1817 = {1{`RANDOM}};
  _T_1267 = _RAND_1817[0:0];
  _RAND_1818 = {1{`RANDOM}};
  _T_1268 = _RAND_1818[0:0];
  _RAND_1819 = {1{`RANDOM}};
  _T_1269 = _RAND_1819[0:0];
  _RAND_1820 = {1{`RANDOM}};
  _T_1270 = _RAND_1820[0:0];
  _RAND_1821 = {1{`RANDOM}};
  _T_1271 = _RAND_1821[0:0];
  _RAND_1822 = {1{`RANDOM}};
  _T_1272 = _RAND_1822[0:0];
  _RAND_1823 = {1{`RANDOM}};
  _T_1273 = _RAND_1823[0:0];
  _RAND_1824 = {1{`RANDOM}};
  _T_1274 = _RAND_1824[0:0];
  _RAND_1825 = {1{`RANDOM}};
  _T_1275 = _RAND_1825[0:0];
  _RAND_1826 = {1{`RANDOM}};
  _T_1276 = _RAND_1826[0:0];
  _RAND_1827 = {1{`RANDOM}};
  _T_1277 = _RAND_1827[0:0];
  _RAND_1828 = {1{`RANDOM}};
  _T_1278 = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  _T_1279 = _RAND_1829[0:0];
  _RAND_1830 = {1{`RANDOM}};
  _T_1280 = _RAND_1830[0:0];
  _RAND_1831 = {1{`RANDOM}};
  _T_1281 = _RAND_1831[0:0];
  _RAND_1832 = {1{`RANDOM}};
  _T_1282 = _RAND_1832[0:0];
  _RAND_1833 = {1{`RANDOM}};
  _T_1283 = _RAND_1833[0:0];
  _RAND_1834 = {1{`RANDOM}};
  _T_1284 = _RAND_1834[0:0];
  _RAND_1835 = {1{`RANDOM}};
  _T_1285 = _RAND_1835[0:0];
  _RAND_1836 = {1{`RANDOM}};
  _T_1286 = _RAND_1836[0:0];
  _RAND_1837 = {1{`RANDOM}};
  _T_1287 = _RAND_1837[0:0];
  _RAND_1838 = {1{`RANDOM}};
  _T_1288 = _RAND_1838[0:0];
  _RAND_1839 = {1{`RANDOM}};
  _T_1289 = _RAND_1839[0:0];
  _RAND_1840 = {1{`RANDOM}};
  _T_1290 = _RAND_1840[0:0];
  _RAND_1841 = {1{`RANDOM}};
  _T_1291 = _RAND_1841[0:0];
  _RAND_1842 = {1{`RANDOM}};
  _T_1292 = _RAND_1842[0:0];
  _RAND_1843 = {1{`RANDOM}};
  _T_1293 = _RAND_1843[0:0];
  _RAND_1844 = {1{`RANDOM}};
  _T_1294 = _RAND_1844[0:0];
  _RAND_1845 = {1{`RANDOM}};
  _T_1295 = _RAND_1845[0:0];
  _RAND_1846 = {1{`RANDOM}};
  _T_1296 = _RAND_1846[0:0];
  _RAND_1847 = {1{`RANDOM}};
  _T_1297 = _RAND_1847[0:0];
  _RAND_1848 = {1{`RANDOM}};
  _T_1298 = _RAND_1848[0:0];
  _RAND_1849 = {1{`RANDOM}};
  _T_1299 = _RAND_1849[0:0];
  _RAND_1850 = {1{`RANDOM}};
  _T_1300 = _RAND_1850[0:0];
  _RAND_1851 = {1{`RANDOM}};
  _T_1301 = _RAND_1851[0:0];
  _RAND_1852 = {1{`RANDOM}};
  _T_1302 = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  _T_1303 = _RAND_1853[0:0];
  _RAND_1854 = {1{`RANDOM}};
  _T_1304 = _RAND_1854[0:0];
  _RAND_1855 = {1{`RANDOM}};
  _T_1305 = _RAND_1855[0:0];
  _RAND_1856 = {1{`RANDOM}};
  _T_1306 = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  _T_1307 = _RAND_1857[0:0];
  _RAND_1858 = {1{`RANDOM}};
  _T_1308 = _RAND_1858[0:0];
  _RAND_1859 = {1{`RANDOM}};
  _T_1309 = _RAND_1859[0:0];
  _RAND_1860 = {1{`RANDOM}};
  _T_1310 = _RAND_1860[0:0];
  _RAND_1861 = {1{`RANDOM}};
  _T_1311 = _RAND_1861[0:0];
  _RAND_1862 = {1{`RANDOM}};
  _T_1312 = _RAND_1862[0:0];
  _RAND_1863 = {1{`RANDOM}};
  _T_1313 = _RAND_1863[0:0];
  _RAND_1864 = {1{`RANDOM}};
  _T_1314 = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  _T_1315 = _RAND_1865[0:0];
  _RAND_1866 = {1{`RANDOM}};
  _T_1316 = _RAND_1866[0:0];
  _RAND_1867 = {1{`RANDOM}};
  _T_1317 = _RAND_1867[0:0];
  _RAND_1868 = {1{`RANDOM}};
  _T_1318 = _RAND_1868[0:0];
  _RAND_1869 = {1{`RANDOM}};
  _T_1319 = _RAND_1869[0:0];
  _RAND_1870 = {1{`RANDOM}};
  _T_1320 = _RAND_1870[0:0];
  _RAND_1871 = {1{`RANDOM}};
  _T_1321 = _RAND_1871[0:0];
  _RAND_1872 = {1{`RANDOM}};
  _T_1322 = _RAND_1872[0:0];
  _RAND_1873 = {1{`RANDOM}};
  _T_1323 = _RAND_1873[0:0];
  _RAND_1874 = {1{`RANDOM}};
  _T_1324 = _RAND_1874[0:0];
  _RAND_1875 = {1{`RANDOM}};
  _T_1325 = _RAND_1875[0:0];
  _RAND_1876 = {1{`RANDOM}};
  _T_1326 = _RAND_1876[0:0];
  _RAND_1877 = {1{`RANDOM}};
  _T_1327 = _RAND_1877[0:0];
  _RAND_1878 = {1{`RANDOM}};
  _T_1328 = _RAND_1878[0:0];
  _RAND_1879 = {1{`RANDOM}};
  _T_1329 = _RAND_1879[0:0];
  _RAND_1880 = {1{`RANDOM}};
  _T_1330 = _RAND_1880[0:0];
  _RAND_1881 = {1{`RANDOM}};
  _T_1331 = _RAND_1881[0:0];
  _RAND_1882 = {1{`RANDOM}};
  _T_1332 = _RAND_1882[0:0];
  _RAND_1883 = {1{`RANDOM}};
  _T_1333 = _RAND_1883[0:0];
  _RAND_1884 = {1{`RANDOM}};
  _T_1334 = _RAND_1884[0:0];
  _RAND_1885 = {1{`RANDOM}};
  _T_1335 = _RAND_1885[0:0];
  _RAND_1886 = {1{`RANDOM}};
  _T_1336 = _RAND_1886[0:0];
  _RAND_1887 = {1{`RANDOM}};
  _T_1337 = _RAND_1887[0:0];
  _RAND_1888 = {1{`RANDOM}};
  _T_1338 = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  _T_1339 = _RAND_1889[0:0];
  _RAND_1890 = {1{`RANDOM}};
  _T_1340 = _RAND_1890[0:0];
  _RAND_1891 = {1{`RANDOM}};
  _T_1341 = _RAND_1891[0:0];
  _RAND_1892 = {1{`RANDOM}};
  _T_1342 = _RAND_1892[0:0];
  _RAND_1893 = {1{`RANDOM}};
  _T_1343 = _RAND_1893[0:0];
  _RAND_1894 = {1{`RANDOM}};
  _T_1344 = _RAND_1894[0:0];
  _RAND_1895 = {1{`RANDOM}};
  _T_1345 = _RAND_1895[0:0];
  _RAND_1896 = {1{`RANDOM}};
  _T_1346 = _RAND_1896[0:0];
  _RAND_1897 = {1{`RANDOM}};
  _T_1347 = _RAND_1897[0:0];
  _RAND_1898 = {1{`RANDOM}};
  _T_1348 = _RAND_1898[0:0];
  _RAND_1899 = {1{`RANDOM}};
  _T_1349 = _RAND_1899[0:0];
  _RAND_1900 = {1{`RANDOM}};
  _T_1350 = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  _T_1351 = _RAND_1901[0:0];
  _RAND_1902 = {1{`RANDOM}};
  _T_1352 = _RAND_1902[0:0];
  _RAND_1903 = {1{`RANDOM}};
  _T_1353 = _RAND_1903[0:0];
  _RAND_1904 = {1{`RANDOM}};
  _T_1354 = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  _T_1355 = _RAND_1905[0:0];
  _RAND_1906 = {1{`RANDOM}};
  _T_1356 = _RAND_1906[0:0];
  _RAND_1907 = {1{`RANDOM}};
  _T_1357 = _RAND_1907[0:0];
  _RAND_1908 = {1{`RANDOM}};
  _T_1358 = _RAND_1908[0:0];
  _RAND_1909 = {1{`RANDOM}};
  _T_1359 = _RAND_1909[0:0];
  _RAND_1910 = {1{`RANDOM}};
  _T_1360 = _RAND_1910[0:0];
  _RAND_1911 = {1{`RANDOM}};
  _T_1361 = _RAND_1911[0:0];
  _RAND_1912 = {1{`RANDOM}};
  _T_1362 = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  _T_1363 = _RAND_1913[0:0];
  _RAND_1914 = {1{`RANDOM}};
  _T_1364 = _RAND_1914[0:0];
  _RAND_1915 = {1{`RANDOM}};
  _T_1365 = _RAND_1915[0:0];
  _RAND_1916 = {1{`RANDOM}};
  _T_1366 = _RAND_1916[0:0];
  _RAND_1917 = {1{`RANDOM}};
  _T_1367 = _RAND_1917[0:0];
  _RAND_1918 = {1{`RANDOM}};
  _T_1368 = _RAND_1918[0:0];
  _RAND_1919 = {1{`RANDOM}};
  _T_1369 = _RAND_1919[0:0];
  _RAND_1920 = {1{`RANDOM}};
  _T_1370 = _RAND_1920[0:0];
  _RAND_1921 = {1{`RANDOM}};
  _T_1371 = _RAND_1921[0:0];
  _RAND_1922 = {1{`RANDOM}};
  _T_1372 = _RAND_1922[0:0];
  _RAND_1923 = {1{`RANDOM}};
  _T_1373 = _RAND_1923[0:0];
  _RAND_1924 = {1{`RANDOM}};
  _T_1374 = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  _T_1375 = _RAND_1925[0:0];
  _RAND_1926 = {1{`RANDOM}};
  _T_1376 = _RAND_1926[0:0];
  _RAND_1927 = {1{`RANDOM}};
  _T_1377 = _RAND_1927[0:0];
  _RAND_1928 = {1{`RANDOM}};
  _T_1378 = _RAND_1928[0:0];
  _RAND_1929 = {1{`RANDOM}};
  _T_1379 = _RAND_1929[0:0];
  _RAND_1930 = {1{`RANDOM}};
  _T_1380 = _RAND_1930[0:0];
  _RAND_1931 = {1{`RANDOM}};
  _T_1381 = _RAND_1931[0:0];
  _RAND_1932 = {1{`RANDOM}};
  _T_1382 = _RAND_1932[0:0];
  _RAND_1933 = {1{`RANDOM}};
  _T_1383 = _RAND_1933[0:0];
  _RAND_1934 = {1{`RANDOM}};
  _T_1384 = _RAND_1934[0:0];
  _RAND_1935 = {1{`RANDOM}};
  _T_1385 = _RAND_1935[0:0];
  _RAND_1936 = {1{`RANDOM}};
  _T_1386 = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  _T_1387 = _RAND_1937[0:0];
  _RAND_1938 = {1{`RANDOM}};
  _T_1388 = _RAND_1938[0:0];
  _RAND_1939 = {1{`RANDOM}};
  _T_1389 = _RAND_1939[0:0];
  _RAND_1940 = {1{`RANDOM}};
  _T_1390 = _RAND_1940[0:0];
  _RAND_1941 = {1{`RANDOM}};
  _T_1391 = _RAND_1941[0:0];
  _RAND_1942 = {1{`RANDOM}};
  _T_1392 = _RAND_1942[0:0];
  _RAND_1943 = {1{`RANDOM}};
  _T_1393 = _RAND_1943[0:0];
  _RAND_1944 = {1{`RANDOM}};
  _T_1394 = _RAND_1944[0:0];
  _RAND_1945 = {1{`RANDOM}};
  _T_1395 = _RAND_1945[0:0];
  _RAND_1946 = {1{`RANDOM}};
  _T_1396 = _RAND_1946[0:0];
  _RAND_1947 = {1{`RANDOM}};
  _T_1397 = _RAND_1947[0:0];
  _RAND_1948 = {1{`RANDOM}};
  _T_1398 = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  _T_1399 = _RAND_1949[0:0];
  _RAND_1950 = {1{`RANDOM}};
  _T_1400 = _RAND_1950[0:0];
  _RAND_1951 = {1{`RANDOM}};
  _T_1401 = _RAND_1951[0:0];
  _RAND_1952 = {1{`RANDOM}};
  _T_1402 = _RAND_1952[0:0];
  _RAND_1953 = {1{`RANDOM}};
  _T_1403 = _RAND_1953[0:0];
  _RAND_1954 = {1{`RANDOM}};
  _T_1404 = _RAND_1954[0:0];
  _RAND_1955 = {1{`RANDOM}};
  _T_1405 = _RAND_1955[0:0];
  _RAND_1956 = {1{`RANDOM}};
  _T_1406 = _RAND_1956[0:0];
  _RAND_1957 = {1{`RANDOM}};
  _T_1407 = _RAND_1957[0:0];
  _RAND_1958 = {1{`RANDOM}};
  _T_1408 = _RAND_1958[0:0];
  _RAND_1959 = {1{`RANDOM}};
  _T_1409 = _RAND_1959[0:0];
  _RAND_1960 = {1{`RANDOM}};
  _T_1410 = _RAND_1960[0:0];
  _RAND_1961 = {1{`RANDOM}};
  _T_1411 = _RAND_1961[0:0];
  _RAND_1962 = {1{`RANDOM}};
  _T_1412 = _RAND_1962[0:0];
  _RAND_1963 = {1{`RANDOM}};
  _T_1413 = _RAND_1963[0:0];
  _RAND_1964 = {1{`RANDOM}};
  _T_1414 = _RAND_1964[0:0];
  _RAND_1965 = {1{`RANDOM}};
  _T_1415 = _RAND_1965[0:0];
  _RAND_1966 = {1{`RANDOM}};
  _T_1416 = _RAND_1966[0:0];
  _RAND_1967 = {1{`RANDOM}};
  _T_1417 = _RAND_1967[0:0];
  _RAND_1968 = {1{`RANDOM}};
  _T_1418 = _RAND_1968[0:0];
  _RAND_1969 = {1{`RANDOM}};
  _T_1419 = _RAND_1969[0:0];
  _RAND_1970 = {1{`RANDOM}};
  _T_1420 = _RAND_1970[0:0];
  _RAND_1971 = {1{`RANDOM}};
  _T_1421 = _RAND_1971[0:0];
  _RAND_1972 = {1{`RANDOM}};
  _T_1422 = _RAND_1972[0:0];
  _RAND_1973 = {1{`RANDOM}};
  _T_1423 = _RAND_1973[0:0];
  _RAND_1974 = {1{`RANDOM}};
  _T_1424 = _RAND_1974[0:0];
  _RAND_1975 = {1{`RANDOM}};
  _T_1425 = _RAND_1975[0:0];
  _RAND_1976 = {1{`RANDOM}};
  _T_1426 = _RAND_1976[0:0];
  _RAND_1977 = {1{`RANDOM}};
  _T_1427 = _RAND_1977[0:0];
  _RAND_1978 = {1{`RANDOM}};
  _T_1428 = _RAND_1978[0:0];
  _RAND_1979 = {1{`RANDOM}};
  _T_1429 = _RAND_1979[0:0];
  _RAND_1980 = {1{`RANDOM}};
  _T_1430 = _RAND_1980[0:0];
  _RAND_1981 = {1{`RANDOM}};
  _T_1431 = _RAND_1981[0:0];
  _RAND_1982 = {1{`RANDOM}};
  _T_1432 = _RAND_1982[0:0];
  _RAND_1983 = {1{`RANDOM}};
  _T_1433 = _RAND_1983[0:0];
  _RAND_1984 = {1{`RANDOM}};
  _T_1434 = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  _T_1435 = _RAND_1985[0:0];
  _RAND_1986 = {1{`RANDOM}};
  _T_1436 = _RAND_1986[0:0];
  _RAND_1987 = {1{`RANDOM}};
  _T_1437 = _RAND_1987[0:0];
  _RAND_1988 = {1{`RANDOM}};
  _T_1438 = _RAND_1988[0:0];
  _RAND_1989 = {1{`RANDOM}};
  _T_1439 = _RAND_1989[0:0];
  _RAND_1990 = {1{`RANDOM}};
  _T_1440 = _RAND_1990[0:0];
  _RAND_1991 = {1{`RANDOM}};
  _T_1441 = _RAND_1991[0:0];
  _RAND_1992 = {1{`RANDOM}};
  _T_1442 = _RAND_1992[0:0];
  _RAND_1993 = {1{`RANDOM}};
  _T_1443 = _RAND_1993[0:0];
  _RAND_1994 = {1{`RANDOM}};
  _T_1444 = _RAND_1994[0:0];
  _RAND_1995 = {1{`RANDOM}};
  _T_1445 = _RAND_1995[0:0];
  _RAND_1996 = {1{`RANDOM}};
  _T_1446 = _RAND_1996[0:0];
  _RAND_1997 = {1{`RANDOM}};
  _T_1447 = _RAND_1997[0:0];
  _RAND_1998 = {1{`RANDOM}};
  _T_1448 = _RAND_1998[0:0];
  _RAND_1999 = {1{`RANDOM}};
  _T_1449 = _RAND_1999[0:0];
  _RAND_2000 = {1{`RANDOM}};
  _T_1450 = _RAND_2000[0:0];
  _RAND_2001 = {1{`RANDOM}};
  _T_1451 = _RAND_2001[0:0];
  _RAND_2002 = {1{`RANDOM}};
  _T_1452 = _RAND_2002[0:0];
  _RAND_2003 = {1{`RANDOM}};
  _T_1453 = _RAND_2003[0:0];
  _RAND_2004 = {1{`RANDOM}};
  _T_1454 = _RAND_2004[0:0];
  _RAND_2005 = {1{`RANDOM}};
  _T_1455 = _RAND_2005[0:0];
  _RAND_2006 = {1{`RANDOM}};
  _T_1456 = _RAND_2006[0:0];
  _RAND_2007 = {1{`RANDOM}};
  _T_1457 = _RAND_2007[0:0];
  _RAND_2008 = {1{`RANDOM}};
  _T_1458 = _RAND_2008[0:0];
  _RAND_2009 = {1{`RANDOM}};
  _T_1459 = _RAND_2009[0:0];
  _RAND_2010 = {1{`RANDOM}};
  _T_1460 = _RAND_2010[0:0];
  _RAND_2011 = {1{`RANDOM}};
  _T_1461 = _RAND_2011[0:0];
  _RAND_2012 = {1{`RANDOM}};
  _T_1462 = _RAND_2012[0:0];
  _RAND_2013 = {1{`RANDOM}};
  _T_1463 = _RAND_2013[0:0];
  _RAND_2014 = {1{`RANDOM}};
  _T_1464 = _RAND_2014[0:0];
  _RAND_2015 = {1{`RANDOM}};
  _T_1465 = _RAND_2015[0:0];
  _RAND_2016 = {1{`RANDOM}};
  _T_1466 = _RAND_2016[0:0];
  _RAND_2017 = {1{`RANDOM}};
  _T_1467 = _RAND_2017[0:0];
  _RAND_2018 = {1{`RANDOM}};
  _T_1468 = _RAND_2018[0:0];
  _RAND_2019 = {1{`RANDOM}};
  _T_1469 = _RAND_2019[0:0];
  _RAND_2020 = {1{`RANDOM}};
  _T_1470 = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  _T_1471 = _RAND_2021[0:0];
  _RAND_2022 = {1{`RANDOM}};
  _T_1472 = _RAND_2022[0:0];
  _RAND_2023 = {1{`RANDOM}};
  _T_1473 = _RAND_2023[0:0];
  _RAND_2024 = {1{`RANDOM}};
  _T_1474 = _RAND_2024[0:0];
  _RAND_2025 = {1{`RANDOM}};
  _T_1475 = _RAND_2025[0:0];
  _RAND_2026 = {1{`RANDOM}};
  _T_1476 = _RAND_2026[0:0];
  _RAND_2027 = {1{`RANDOM}};
  _T_1477 = _RAND_2027[0:0];
  _RAND_2028 = {1{`RANDOM}};
  _T_1478 = _RAND_2028[0:0];
  _RAND_2029 = {1{`RANDOM}};
  _T_1479 = _RAND_2029[0:0];
  _RAND_2030 = {1{`RANDOM}};
  _T_1480 = _RAND_2030[0:0];
  _RAND_2031 = {1{`RANDOM}};
  _T_1481 = _RAND_2031[0:0];
  _RAND_2032 = {1{`RANDOM}};
  _T_1482 = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  _T_1483 = _RAND_2033[0:0];
  _RAND_2034 = {1{`RANDOM}};
  _T_1484 = _RAND_2034[0:0];
  _RAND_2035 = {1{`RANDOM}};
  _T_1485 = _RAND_2035[0:0];
  _RAND_2036 = {1{`RANDOM}};
  _T_1486 = _RAND_2036[0:0];
  _RAND_2037 = {1{`RANDOM}};
  _T_1487 = _RAND_2037[0:0];
  _RAND_2038 = {1{`RANDOM}};
  _T_1488 = _RAND_2038[0:0];
  _RAND_2039 = {1{`RANDOM}};
  _T_1489 = _RAND_2039[0:0];
  _RAND_2040 = {1{`RANDOM}};
  _T_1490 = _RAND_2040[0:0];
  _RAND_2041 = {1{`RANDOM}};
  _T_1491 = _RAND_2041[0:0];
  _RAND_2042 = {1{`RANDOM}};
  _T_1492 = _RAND_2042[0:0];
  _RAND_2043 = {1{`RANDOM}};
  _T_1493 = _RAND_2043[0:0];
  _RAND_2044 = {1{`RANDOM}};
  _T_1494 = _RAND_2044[0:0];
  _RAND_2045 = {1{`RANDOM}};
  _T_1495 = _RAND_2045[0:0];
  _RAND_2046 = {1{`RANDOM}};
  _T_1496 = _RAND_2046[0:0];
  _RAND_2047 = {1{`RANDOM}};
  _T_1497 = _RAND_2047[0:0];
  _RAND_2048 = {1{`RANDOM}};
  _T_1498 = _RAND_2048[0:0];
  _RAND_2049 = {1{`RANDOM}};
  _T_1499 = _RAND_2049[0:0];
  _RAND_2050 = {1{`RANDOM}};
  _T_1500 = _RAND_2050[0:0];
  _RAND_2051 = {1{`RANDOM}};
  _T_1501 = _RAND_2051[0:0];
  _RAND_2052 = {1{`RANDOM}};
  _T_1502 = _RAND_2052[0:0];
  _RAND_2053 = {1{`RANDOM}};
  _T_1503 = _RAND_2053[0:0];
  _RAND_2054 = {1{`RANDOM}};
  _T_1504 = _RAND_2054[0:0];
  _RAND_2055 = {1{`RANDOM}};
  _T_1505 = _RAND_2055[0:0];
  _RAND_2056 = {1{`RANDOM}};
  _T_1506 = _RAND_2056[0:0];
  _RAND_2057 = {1{`RANDOM}};
  _T_1507 = _RAND_2057[0:0];
  _RAND_2058 = {1{`RANDOM}};
  _T_1508 = _RAND_2058[0:0];
  _RAND_2059 = {1{`RANDOM}};
  _T_1509 = _RAND_2059[0:0];
  _RAND_2060 = {1{`RANDOM}};
  _T_1510 = _RAND_2060[0:0];
  _RAND_2061 = {1{`RANDOM}};
  _T_1511 = _RAND_2061[0:0];
  _RAND_2062 = {1{`RANDOM}};
  _T_1512 = _RAND_2062[0:0];
  _RAND_2063 = {1{`RANDOM}};
  _T_1513 = _RAND_2063[0:0];
  _RAND_2064 = {1{`RANDOM}};
  _T_1514 = _RAND_2064[0:0];
  _RAND_2065 = {1{`RANDOM}};
  _T_1515 = _RAND_2065[0:0];
  _RAND_2066 = {1{`RANDOM}};
  _T_1516 = _RAND_2066[0:0];
  _RAND_2067 = {1{`RANDOM}};
  _T_1517 = _RAND_2067[0:0];
  _RAND_2068 = {1{`RANDOM}};
  _T_1518 = _RAND_2068[0:0];
  _RAND_2069 = {1{`RANDOM}};
  _T_1519 = _RAND_2069[0:0];
  _RAND_2070 = {1{`RANDOM}};
  _T_1520 = _RAND_2070[0:0];
  _RAND_2071 = {1{`RANDOM}};
  _T_1521 = _RAND_2071[0:0];
  _RAND_2072 = {1{`RANDOM}};
  _T_1522 = _RAND_2072[0:0];
  _RAND_2073 = {1{`RANDOM}};
  _T_1523 = _RAND_2073[0:0];
  _RAND_2074 = {1{`RANDOM}};
  _T_1524 = _RAND_2074[0:0];
  _RAND_2075 = {1{`RANDOM}};
  _T_1525 = _RAND_2075[0:0];
  _RAND_2076 = {1{`RANDOM}};
  _T_1526 = _RAND_2076[0:0];
  _RAND_2077 = {1{`RANDOM}};
  _T_1527 = _RAND_2077[0:0];
  _RAND_2078 = {1{`RANDOM}};
  _T_1528 = _RAND_2078[0:0];
  _RAND_2079 = {1{`RANDOM}};
  _T_1529 = _RAND_2079[0:0];
  _RAND_2080 = {1{`RANDOM}};
  _T_1530 = _RAND_2080[0:0];
  _RAND_2081 = {1{`RANDOM}};
  _T_1531 = _RAND_2081[0:0];
  _RAND_2082 = {1{`RANDOM}};
  _T_1532 = _RAND_2082[0:0];
  _RAND_2083 = {1{`RANDOM}};
  _T_1533 = _RAND_2083[0:0];
  _RAND_2084 = {1{`RANDOM}};
  _T_1534 = _RAND_2084[0:0];
  _RAND_2085 = {1{`RANDOM}};
  _T_1535 = _RAND_2085[0:0];
  _RAND_2086 = {1{`RANDOM}};
  _T_1536 = _RAND_2086[0:0];
  _RAND_2087 = {1{`RANDOM}};
  _T_1537 = _RAND_2087[0:0];
  _RAND_2088 = {1{`RANDOM}};
  _T_1538 = _RAND_2088[0:0];
  _RAND_2089 = {1{`RANDOM}};
  _T_1539 = _RAND_2089[0:0];
  _RAND_2090 = {1{`RANDOM}};
  _T_1540 = _RAND_2090[0:0];
  _RAND_2091 = {1{`RANDOM}};
  _T_1541 = _RAND_2091[0:0];
  _RAND_2092 = {1{`RANDOM}};
  _T_1542 = _RAND_2092[0:0];
  _RAND_2093 = {1{`RANDOM}};
  _T_1543 = _RAND_2093[0:0];
  _RAND_2094 = {1{`RANDOM}};
  _T_1544 = _RAND_2094[0:0];
  _RAND_2095 = {1{`RANDOM}};
  _T_1545 = _RAND_2095[0:0];
  _RAND_2096 = {1{`RANDOM}};
  _T_1546 = _RAND_2096[0:0];
  _RAND_2097 = {1{`RANDOM}};
  _T_1547 = _RAND_2097[0:0];
  _RAND_2098 = {1{`RANDOM}};
  _T_1548 = _RAND_2098[0:0];
  _RAND_2099 = {1{`RANDOM}};
  _T_1549 = _RAND_2099[0:0];
  _RAND_2100 = {1{`RANDOM}};
  _T_1550 = _RAND_2100[0:0];
  _RAND_2101 = {1{`RANDOM}};
  _T_1551 = _RAND_2101[0:0];
  _RAND_2102 = {1{`RANDOM}};
  _T_1552 = _RAND_2102[0:0];
  _RAND_2103 = {1{`RANDOM}};
  _T_1553 = _RAND_2103[0:0];
  _RAND_2104 = {1{`RANDOM}};
  _T_1554 = _RAND_2104[0:0];
  _RAND_2105 = {1{`RANDOM}};
  _T_1555 = _RAND_2105[0:0];
  _RAND_2106 = {1{`RANDOM}};
  _T_1556 = _RAND_2106[0:0];
  _RAND_2107 = {1{`RANDOM}};
  _T_1557 = _RAND_2107[0:0];
  _RAND_2108 = {1{`RANDOM}};
  _T_1558 = _RAND_2108[0:0];
  _RAND_2109 = {1{`RANDOM}};
  _T_1559 = _RAND_2109[0:0];
  _RAND_2110 = {1{`RANDOM}};
  _T_1560 = _RAND_2110[0:0];
  _RAND_2111 = {1{`RANDOM}};
  _T_1561 = _RAND_2111[0:0];
  _RAND_2112 = {1{`RANDOM}};
  _T_1562 = _RAND_2112[0:0];
  _RAND_2113 = {1{`RANDOM}};
  _T_1563 = _RAND_2113[0:0];
  _RAND_2114 = {1{`RANDOM}};
  _T_1564 = _RAND_2114[0:0];
  _RAND_2115 = {1{`RANDOM}};
  _T_1565 = _RAND_2115[0:0];
  _RAND_2116 = {1{`RANDOM}};
  _T_1566 = _RAND_2116[0:0];
  _RAND_2117 = {1{`RANDOM}};
  _T_1567 = _RAND_2117[0:0];
  _RAND_2118 = {1{`RANDOM}};
  _T_1568 = _RAND_2118[0:0];
  _RAND_2119 = {1{`RANDOM}};
  _T_1569 = _RAND_2119[0:0];
  _RAND_2120 = {1{`RANDOM}};
  _T_1570 = _RAND_2120[0:0];
  _RAND_2121 = {1{`RANDOM}};
  _T_1571 = _RAND_2121[0:0];
  _RAND_2122 = {1{`RANDOM}};
  _T_1572 = _RAND_2122[0:0];
  _RAND_2123 = {1{`RANDOM}};
  _T_1573 = _RAND_2123[0:0];
  _RAND_2124 = {1{`RANDOM}};
  _T_1574 = _RAND_2124[0:0];
  _RAND_2125 = {1{`RANDOM}};
  _T_1575 = _RAND_2125[0:0];
  _RAND_2126 = {1{`RANDOM}};
  _T_1576 = _RAND_2126[0:0];
  _RAND_2127 = {1{`RANDOM}};
  _T_1577 = _RAND_2127[0:0];
  _RAND_2128 = {1{`RANDOM}};
  _T_1578 = _RAND_2128[0:0];
  _RAND_2129 = {1{`RANDOM}};
  _T_1579 = _RAND_2129[0:0];
  _RAND_2130 = {1{`RANDOM}};
  _T_1580 = _RAND_2130[0:0];
  _RAND_2131 = {1{`RANDOM}};
  _T_1581 = _RAND_2131[0:0];
  _RAND_2132 = {1{`RANDOM}};
  _T_1582 = _RAND_2132[0:0];
  _RAND_2133 = {1{`RANDOM}};
  _T_1583 = _RAND_2133[0:0];
  _RAND_2134 = {1{`RANDOM}};
  _T_1584 = _RAND_2134[0:0];
  _RAND_2135 = {1{`RANDOM}};
  _T_1585 = _RAND_2135[0:0];
  _RAND_2136 = {1{`RANDOM}};
  _T_1586 = _RAND_2136[0:0];
  _RAND_2137 = {1{`RANDOM}};
  _T_1587 = _RAND_2137[0:0];
  _RAND_2138 = {1{`RANDOM}};
  _T_1588 = _RAND_2138[0:0];
  _RAND_2139 = {1{`RANDOM}};
  _T_1589 = _RAND_2139[0:0];
  _RAND_2140 = {1{`RANDOM}};
  _T_1590 = _RAND_2140[0:0];
  _RAND_2141 = {1{`RANDOM}};
  _T_1591 = _RAND_2141[0:0];
  _RAND_2142 = {1{`RANDOM}};
  _T_1592 = _RAND_2142[0:0];
  _RAND_2143 = {1{`RANDOM}};
  _T_1593 = _RAND_2143[0:0];
  _RAND_2144 = {1{`RANDOM}};
  _T_1594 = _RAND_2144[0:0];
  _RAND_2145 = {1{`RANDOM}};
  _T_1595 = _RAND_2145[0:0];
  _RAND_2146 = {1{`RANDOM}};
  _T_1596 = _RAND_2146[0:0];
  _RAND_2147 = {1{`RANDOM}};
  _T_1597 = _RAND_2147[0:0];
  _RAND_2148 = {1{`RANDOM}};
  _T_1598 = _RAND_2148[0:0];
  _RAND_2149 = {1{`RANDOM}};
  _T_1599 = _RAND_2149[0:0];
  _RAND_2150 = {1{`RANDOM}};
  _T_1600 = _RAND_2150[0:0];
  _RAND_2151 = {1{`RANDOM}};
  _T_1601 = _RAND_2151[0:0];
  _RAND_2152 = {1{`RANDOM}};
  _T_1602 = _RAND_2152[0:0];
  _RAND_2153 = {1{`RANDOM}};
  _T_1603 = _RAND_2153[0:0];
  _RAND_2154 = {1{`RANDOM}};
  _T_1604 = _RAND_2154[0:0];
  _RAND_2155 = {1{`RANDOM}};
  _T_1605 = _RAND_2155[0:0];
  _RAND_2156 = {1{`RANDOM}};
  _T_1606 = _RAND_2156[0:0];
  _RAND_2157 = {1{`RANDOM}};
  _T_1607 = _RAND_2157[0:0];
  _RAND_2158 = {1{`RANDOM}};
  _T_1608 = _RAND_2158[0:0];
  _RAND_2159 = {1{`RANDOM}};
  _T_1609 = _RAND_2159[0:0];
  _RAND_2160 = {1{`RANDOM}};
  _T_1610 = _RAND_2160[0:0];
  _RAND_2161 = {1{`RANDOM}};
  _T_1611 = _RAND_2161[0:0];
  _RAND_2162 = {1{`RANDOM}};
  _T_1612 = _RAND_2162[0:0];
  _RAND_2163 = {1{`RANDOM}};
  _T_1613 = _RAND_2163[0:0];
  _RAND_2164 = {1{`RANDOM}};
  _T_1614 = _RAND_2164[0:0];
  _RAND_2165 = {1{`RANDOM}};
  _T_1615 = _RAND_2165[0:0];
  _RAND_2166 = {1{`RANDOM}};
  _T_1616 = _RAND_2166[0:0];
  _RAND_2167 = {1{`RANDOM}};
  _T_1617 = _RAND_2167[0:0];
  _RAND_2168 = {1{`RANDOM}};
  _T_1618 = _RAND_2168[0:0];
  _RAND_2169 = {1{`RANDOM}};
  _T_1619 = _RAND_2169[0:0];
  _RAND_2170 = {1{`RANDOM}};
  _T_1620 = _RAND_2170[0:0];
  _RAND_2171 = {1{`RANDOM}};
  _T_1621 = _RAND_2171[0:0];
  _RAND_2172 = {1{`RANDOM}};
  _T_1622 = _RAND_2172[0:0];
  _RAND_2173 = {1{`RANDOM}};
  _T_1623 = _RAND_2173[0:0];
  _RAND_2174 = {1{`RANDOM}};
  _T_1624 = _RAND_2174[0:0];
  _RAND_2175 = {1{`RANDOM}};
  _T_1625 = _RAND_2175[0:0];
  _RAND_2176 = {1{`RANDOM}};
  _T_1626 = _RAND_2176[0:0];
  _RAND_2177 = {1{`RANDOM}};
  _T_1627 = _RAND_2177[0:0];
  _RAND_2178 = {1{`RANDOM}};
  _T_1628 = _RAND_2178[0:0];
  _RAND_2179 = {1{`RANDOM}};
  _T_1629 = _RAND_2179[0:0];
  _RAND_2180 = {1{`RANDOM}};
  _T_1630 = _RAND_2180[0:0];
  _RAND_2181 = {1{`RANDOM}};
  _T_1631 = _RAND_2181[0:0];
  _RAND_2182 = {1{`RANDOM}};
  _T_1632 = _RAND_2182[0:0];
  _RAND_2183 = {1{`RANDOM}};
  _T_1633 = _RAND_2183[0:0];
  _RAND_2184 = {1{`RANDOM}};
  _T_1634 = _RAND_2184[0:0];
  _RAND_2185 = {1{`RANDOM}};
  _T_1635 = _RAND_2185[0:0];
  _RAND_2186 = {1{`RANDOM}};
  _T_1636 = _RAND_2186[0:0];
  _RAND_2187 = {1{`RANDOM}};
  _T_1637 = _RAND_2187[0:0];
  _RAND_2188 = {1{`RANDOM}};
  _T_1638 = _RAND_2188[0:0];
  _RAND_2189 = {1{`RANDOM}};
  _T_1639 = _RAND_2189[0:0];
  _RAND_2190 = {1{`RANDOM}};
  _T_1640 = _RAND_2190[0:0];
  _RAND_2191 = {1{`RANDOM}};
  _T_1641 = _RAND_2191[0:0];
  _RAND_2192 = {1{`RANDOM}};
  _T_1642 = _RAND_2192[0:0];
  _RAND_2193 = {1{`RANDOM}};
  _T_1643 = _RAND_2193[0:0];
  _RAND_2194 = {1{`RANDOM}};
  _T_1644 = _RAND_2194[0:0];
  _RAND_2195 = {1{`RANDOM}};
  _T_1645 = _RAND_2195[0:0];
  _RAND_2196 = {1{`RANDOM}};
  _T_1646 = _RAND_2196[0:0];
  _RAND_2197 = {1{`RANDOM}};
  _T_1647 = _RAND_2197[0:0];
  _RAND_2198 = {1{`RANDOM}};
  _T_1648 = _RAND_2198[0:0];
  _RAND_2199 = {1{`RANDOM}};
  _T_1649 = _RAND_2199[0:0];
  _RAND_2200 = {1{`RANDOM}};
  _T_1650 = _RAND_2200[0:0];
  _RAND_2201 = {1{`RANDOM}};
  _T_1651 = _RAND_2201[0:0];
  _RAND_2202 = {1{`RANDOM}};
  _T_1652 = _RAND_2202[0:0];
  _RAND_2203 = {1{`RANDOM}};
  _T_1653 = _RAND_2203[0:0];
  _RAND_2204 = {1{`RANDOM}};
  _T_1654 = _RAND_2204[0:0];
  _RAND_2205 = {1{`RANDOM}};
  _T_1655 = _RAND_2205[0:0];
  _RAND_2206 = {1{`RANDOM}};
  _T_1656 = _RAND_2206[0:0];
  _RAND_2207 = {1{`RANDOM}};
  _T_1657 = _RAND_2207[0:0];
  _RAND_2208 = {1{`RANDOM}};
  _T_1658 = _RAND_2208[0:0];
  _RAND_2209 = {1{`RANDOM}};
  _T_1659 = _RAND_2209[0:0];
  _RAND_2210 = {1{`RANDOM}};
  _T_1660 = _RAND_2210[0:0];
  _RAND_2211 = {1{`RANDOM}};
  _T_1661 = _RAND_2211[0:0];
  _RAND_2212 = {1{`RANDOM}};
  _T_1662 = _RAND_2212[0:0];
  _RAND_2213 = {1{`RANDOM}};
  _T_1663 = _RAND_2213[0:0];
  _RAND_2214 = {1{`RANDOM}};
  _T_1664 = _RAND_2214[0:0];
  _RAND_2215 = {1{`RANDOM}};
  _T_1665 = _RAND_2215[0:0];
  _RAND_2216 = {1{`RANDOM}};
  _T_1666 = _RAND_2216[0:0];
  _RAND_2217 = {1{`RANDOM}};
  _T_1667 = _RAND_2217[0:0];
  _RAND_2218 = {1{`RANDOM}};
  _T_1668 = _RAND_2218[0:0];
  _RAND_2219 = {1{`RANDOM}};
  _T_1669 = _RAND_2219[0:0];
  _RAND_2220 = {1{`RANDOM}};
  _T_1670 = _RAND_2220[0:0];
  _RAND_2221 = {1{`RANDOM}};
  _T_1671 = _RAND_2221[0:0];
  _RAND_2222 = {1{`RANDOM}};
  _T_1672 = _RAND_2222[0:0];
  _RAND_2223 = {1{`RANDOM}};
  _T_1673 = _RAND_2223[0:0];
  _RAND_2224 = {1{`RANDOM}};
  _T_1674 = _RAND_2224[0:0];
  _RAND_2225 = {1{`RANDOM}};
  _T_1675 = _RAND_2225[0:0];
  _RAND_2226 = {1{`RANDOM}};
  _T_1676 = _RAND_2226[0:0];
  _RAND_2227 = {1{`RANDOM}};
  _T_1677 = _RAND_2227[0:0];
  _RAND_2228 = {1{`RANDOM}};
  _T_1678 = _RAND_2228[0:0];
  _RAND_2229 = {1{`RANDOM}};
  _T_1679 = _RAND_2229[0:0];
  _RAND_2230 = {1{`RANDOM}};
  _T_1680 = _RAND_2230[0:0];
  _RAND_2231 = {1{`RANDOM}};
  _T_1681 = _RAND_2231[0:0];
  _RAND_2232 = {1{`RANDOM}};
  _T_1682 = _RAND_2232[0:0];
  _RAND_2233 = {1{`RANDOM}};
  _T_1683 = _RAND_2233[0:0];
  _RAND_2234 = {1{`RANDOM}};
  _T_1684 = _RAND_2234[0:0];
  _RAND_2235 = {1{`RANDOM}};
  _T_1685 = _RAND_2235[0:0];
  _RAND_2236 = {1{`RANDOM}};
  _T_1686 = _RAND_2236[0:0];
  _RAND_2237 = {1{`RANDOM}};
  _T_1687 = _RAND_2237[0:0];
  _RAND_2238 = {1{`RANDOM}};
  _T_1688 = _RAND_2238[0:0];
  _RAND_2239 = {1{`RANDOM}};
  _T_1689 = _RAND_2239[0:0];
  _RAND_2240 = {1{`RANDOM}};
  _T_1690 = _RAND_2240[0:0];
  _RAND_2241 = {1{`RANDOM}};
  _T_1691 = _RAND_2241[0:0];
  _RAND_2242 = {1{`RANDOM}};
  _T_1692 = _RAND_2242[0:0];
  _RAND_2243 = {1{`RANDOM}};
  _T_1693 = _RAND_2243[0:0];
  _RAND_2244 = {1{`RANDOM}};
  _T_1694 = _RAND_2244[0:0];
  _RAND_2245 = {1{`RANDOM}};
  _T_1695 = _RAND_2245[0:0];
  _RAND_2246 = {1{`RANDOM}};
  _T_1696 = _RAND_2246[0:0];
  _RAND_2247 = {1{`RANDOM}};
  _T_1697 = _RAND_2247[0:0];
  _RAND_2248 = {1{`RANDOM}};
  _T_1698 = _RAND_2248[0:0];
  _RAND_2249 = {1{`RANDOM}};
  _T_1699 = _RAND_2249[0:0];
  _RAND_2250 = {1{`RANDOM}};
  _T_1700 = _RAND_2250[0:0];
  _RAND_2251 = {1{`RANDOM}};
  _T_1701 = _RAND_2251[0:0];
  _RAND_2252 = {1{`RANDOM}};
  _T_1702 = _RAND_2252[0:0];
  _RAND_2253 = {1{`RANDOM}};
  _T_1703 = _RAND_2253[0:0];
  _RAND_2254 = {1{`RANDOM}};
  _T_1704 = _RAND_2254[0:0];
  _RAND_2255 = {1{`RANDOM}};
  _T_1705 = _RAND_2255[0:0];
  _RAND_2256 = {1{`RANDOM}};
  _T_1706 = _RAND_2256[0:0];
  _RAND_2257 = {1{`RANDOM}};
  _T_1707 = _RAND_2257[0:0];
  _RAND_2258 = {1{`RANDOM}};
  _T_1708 = _RAND_2258[0:0];
  _RAND_2259 = {1{`RANDOM}};
  _T_1709 = _RAND_2259[0:0];
  _RAND_2260 = {1{`RANDOM}};
  _T_1710 = _RAND_2260[0:0];
  _RAND_2261 = {1{`RANDOM}};
  _T_1711 = _RAND_2261[0:0];
  _RAND_2262 = {1{`RANDOM}};
  _T_1712 = _RAND_2262[0:0];
  _RAND_2263 = {1{`RANDOM}};
  _T_1713 = _RAND_2263[0:0];
  _RAND_2264 = {1{`RANDOM}};
  _T_1714 = _RAND_2264[0:0];
  _RAND_2265 = {1{`RANDOM}};
  _T_1715 = _RAND_2265[0:0];
  _RAND_2266 = {1{`RANDOM}};
  _T_1716 = _RAND_2266[0:0];
  _RAND_2267 = {1{`RANDOM}};
  _T_1717 = _RAND_2267[0:0];
  _RAND_2268 = {1{`RANDOM}};
  _T_1718 = _RAND_2268[0:0];
  _RAND_2269 = {1{`RANDOM}};
  _T_1719 = _RAND_2269[0:0];
  _RAND_2270 = {1{`RANDOM}};
  _T_1720 = _RAND_2270[0:0];
  _RAND_2271 = {1{`RANDOM}};
  _T_1721 = _RAND_2271[0:0];
  _RAND_2272 = {1{`RANDOM}};
  _T_1722 = _RAND_2272[0:0];
  _RAND_2273 = {1{`RANDOM}};
  _T_1723 = _RAND_2273[0:0];
  _RAND_2274 = {1{`RANDOM}};
  _T_1724 = _RAND_2274[0:0];
  _RAND_2275 = {1{`RANDOM}};
  _T_1725 = _RAND_2275[0:0];
  _RAND_2276 = {1{`RANDOM}};
  _T_1726 = _RAND_2276[0:0];
  _RAND_2277 = {1{`RANDOM}};
  _T_1727 = _RAND_2277[0:0];
  _RAND_2278 = {1{`RANDOM}};
  _T_1728 = _RAND_2278[0:0];
  _RAND_2279 = {1{`RANDOM}};
  _T_1729 = _RAND_2279[0:0];
  _RAND_2280 = {1{`RANDOM}};
  _T_1730 = _RAND_2280[0:0];
  _RAND_2281 = {1{`RANDOM}};
  _T_1731 = _RAND_2281[0:0];
  _RAND_2282 = {1{`RANDOM}};
  _T_1732 = _RAND_2282[0:0];
  _RAND_2283 = {1{`RANDOM}};
  _T_1733 = _RAND_2283[0:0];
  _RAND_2284 = {1{`RANDOM}};
  _T_1734 = _RAND_2284[0:0];
  _RAND_2285 = {1{`RANDOM}};
  _T_1735 = _RAND_2285[0:0];
  _RAND_2286 = {1{`RANDOM}};
  _T_1736 = _RAND_2286[0:0];
  _RAND_2287 = {1{`RANDOM}};
  _T_1737 = _RAND_2287[0:0];
  _RAND_2288 = {1{`RANDOM}};
  _T_1738 = _RAND_2288[0:0];
  _RAND_2289 = {1{`RANDOM}};
  _T_1739 = _RAND_2289[0:0];
  _RAND_2290 = {1{`RANDOM}};
  _T_1740 = _RAND_2290[0:0];
  _RAND_2291 = {1{`RANDOM}};
  _T_1741 = _RAND_2291[0:0];
  _RAND_2292 = {1{`RANDOM}};
  _T_1742 = _RAND_2292[0:0];
  _RAND_2293 = {1{`RANDOM}};
  _T_1743 = _RAND_2293[0:0];
  _RAND_2294 = {1{`RANDOM}};
  _T_1744 = _RAND_2294[0:0];
  _RAND_2295 = {1{`RANDOM}};
  _T_1745 = _RAND_2295[0:0];
  _RAND_2296 = {1{`RANDOM}};
  _T_1746 = _RAND_2296[0:0];
  _RAND_2297 = {1{`RANDOM}};
  _T_1747 = _RAND_2297[0:0];
  _RAND_2298 = {1{`RANDOM}};
  _T_1748 = _RAND_2298[0:0];
  _RAND_2299 = {1{`RANDOM}};
  _T_1749 = _RAND_2299[0:0];
  _RAND_2300 = {1{`RANDOM}};
  _T_1750 = _RAND_2300[0:0];
  _RAND_2301 = {1{`RANDOM}};
  _T_1751 = _RAND_2301[0:0];
  _RAND_2302 = {1{`RANDOM}};
  _T_1752 = _RAND_2302[0:0];
  _RAND_2303 = {1{`RANDOM}};
  _T_1753 = _RAND_2303[0:0];
  _RAND_2304 = {1{`RANDOM}};
  _T_1754 = _RAND_2304[0:0];
  _RAND_2305 = {1{`RANDOM}};
  _T_1755 = _RAND_2305[0:0];
  _RAND_2306 = {1{`RANDOM}};
  _T_1756 = _RAND_2306[0:0];
  _RAND_2307 = {1{`RANDOM}};
  _T_1757 = _RAND_2307[0:0];
  _RAND_2308 = {1{`RANDOM}};
  _T_1758 = _RAND_2308[0:0];
  _RAND_2309 = {1{`RANDOM}};
  _T_1759 = _RAND_2309[0:0];
  _RAND_2310 = {1{`RANDOM}};
  _T_1760 = _RAND_2310[0:0];
  _RAND_2311 = {1{`RANDOM}};
  _T_1761 = _RAND_2311[0:0];
  _RAND_2312 = {1{`RANDOM}};
  _T_1762 = _RAND_2312[0:0];
  _RAND_2313 = {1{`RANDOM}};
  _T_1763 = _RAND_2313[0:0];
  _RAND_2314 = {1{`RANDOM}};
  _T_1764 = _RAND_2314[0:0];
  _RAND_2315 = {1{`RANDOM}};
  _T_1765 = _RAND_2315[0:0];
  _RAND_2316 = {1{`RANDOM}};
  _T_1766 = _RAND_2316[0:0];
  _RAND_2317 = {1{`RANDOM}};
  _T_1767 = _RAND_2317[0:0];
  _RAND_2318 = {1{`RANDOM}};
  _T_1768 = _RAND_2318[0:0];
  _RAND_2319 = {1{`RANDOM}};
  _T_1769 = _RAND_2319[0:0];
  _RAND_2320 = {1{`RANDOM}};
  _T_1770 = _RAND_2320[0:0];
  _RAND_2321 = {1{`RANDOM}};
  _T_1771 = _RAND_2321[0:0];
  _RAND_2322 = {1{`RANDOM}};
  _T_1772 = _RAND_2322[0:0];
  _RAND_2323 = {1{`RANDOM}};
  _T_1773 = _RAND_2323[0:0];
  _RAND_2324 = {1{`RANDOM}};
  _T_1774 = _RAND_2324[0:0];
  _RAND_2325 = {1{`RANDOM}};
  _T_1775 = _RAND_2325[0:0];
  _RAND_2326 = {1{`RANDOM}};
  _T_1776 = _RAND_2326[0:0];
  _RAND_2327 = {1{`RANDOM}};
  _T_1777 = _RAND_2327[0:0];
  _RAND_2328 = {1{`RANDOM}};
  _T_1778 = _RAND_2328[0:0];
  _RAND_2329 = {1{`RANDOM}};
  _T_1779 = _RAND_2329[0:0];
  _RAND_2330 = {1{`RANDOM}};
  _T_1780 = _RAND_2330[0:0];
  _RAND_2331 = {1{`RANDOM}};
  _T_1781 = _RAND_2331[0:0];
  _RAND_2332 = {1{`RANDOM}};
  _T_1782 = _RAND_2332[0:0];
  _RAND_2333 = {1{`RANDOM}};
  _T_1783 = _RAND_2333[0:0];
  _RAND_2334 = {1{`RANDOM}};
  _T_1784 = _RAND_2334[0:0];
  _RAND_2335 = {1{`RANDOM}};
  _T_1785 = _RAND_2335[0:0];
  _RAND_2336 = {1{`RANDOM}};
  _T_1786 = _RAND_2336[0:0];
  _RAND_2337 = {1{`RANDOM}};
  _T_1787 = _RAND_2337[0:0];
  _RAND_2338 = {1{`RANDOM}};
  _T_1788 = _RAND_2338[0:0];
  _RAND_2339 = {1{`RANDOM}};
  _T_1789 = _RAND_2339[0:0];
  _RAND_2340 = {1{`RANDOM}};
  _T_1790 = _RAND_2340[0:0];
  _RAND_2341 = {1{`RANDOM}};
  _T_1791 = _RAND_2341[0:0];
  _RAND_2342 = {1{`RANDOM}};
  _T_1792 = _RAND_2342[0:0];
  _RAND_2343 = {1{`RANDOM}};
  _T_1793 = _RAND_2343[0:0];
  _RAND_2344 = {1{`RANDOM}};
  _T_1794 = _RAND_2344[0:0];
  _RAND_2345 = {1{`RANDOM}};
  _T_1795 = _RAND_2345[0:0];
  _RAND_2346 = {1{`RANDOM}};
  _T_1796 = _RAND_2346[0:0];
  _RAND_2347 = {1{`RANDOM}};
  _T_1797 = _RAND_2347[0:0];
  _RAND_2348 = {1{`RANDOM}};
  _T_1798 = _RAND_2348[0:0];
  _RAND_2349 = {1{`RANDOM}};
  _T_1799 = _RAND_2349[0:0];
  _RAND_2350 = {1{`RANDOM}};
  _T_1800 = _RAND_2350[0:0];
  _RAND_2351 = {1{`RANDOM}};
  _T_1801 = _RAND_2351[0:0];
  _RAND_2352 = {1{`RANDOM}};
  _T_1802 = _RAND_2352[0:0];
  _RAND_2353 = {1{`RANDOM}};
  _T_1803 = _RAND_2353[0:0];
  _RAND_2354 = {1{`RANDOM}};
  _T_1804 = _RAND_2354[0:0];
  _RAND_2355 = {1{`RANDOM}};
  _T_1805 = _RAND_2355[0:0];
  _RAND_2356 = {1{`RANDOM}};
  _T_1806 = _RAND_2356[0:0];
  _RAND_2357 = {1{`RANDOM}};
  _T_1807 = _RAND_2357[0:0];
  _RAND_2358 = {1{`RANDOM}};
  _T_1808 = _RAND_2358[0:0];
  _RAND_2359 = {1{`RANDOM}};
  _T_1809 = _RAND_2359[0:0];
  _RAND_2360 = {1{`RANDOM}};
  _T_1810 = _RAND_2360[0:0];
  _RAND_2361 = {1{`RANDOM}};
  _T_1811 = _RAND_2361[0:0];
  _RAND_2362 = {1{`RANDOM}};
  _T_1812 = _RAND_2362[0:0];
  _RAND_2363 = {1{`RANDOM}};
  _T_1813 = _RAND_2363[0:0];
  _RAND_2364 = {1{`RANDOM}};
  _T_1814 = _RAND_2364[0:0];
  _RAND_2365 = {1{`RANDOM}};
  _T_1815 = _RAND_2365[0:0];
  _RAND_2366 = {1{`RANDOM}};
  _T_1816 = _RAND_2366[0:0];
  _RAND_2367 = {1{`RANDOM}};
  _T_1817 = _RAND_2367[0:0];
  _RAND_2368 = {1{`RANDOM}};
  _T_1818 = _RAND_2368[0:0];
  _RAND_2369 = {1{`RANDOM}};
  _T_1819 = _RAND_2369[0:0];
  _RAND_2370 = {1{`RANDOM}};
  _T_1820 = _RAND_2370[0:0];
  _RAND_2371 = {1{`RANDOM}};
  _T_1821 = _RAND_2371[0:0];
  _RAND_2372 = {1{`RANDOM}};
  _T_1822 = _RAND_2372[0:0];
  _RAND_2373 = {1{`RANDOM}};
  _T_1823 = _RAND_2373[0:0];
  _RAND_2374 = {1{`RANDOM}};
  _T_1824 = _RAND_2374[0:0];
  _RAND_2375 = {1{`RANDOM}};
  _T_1825 = _RAND_2375[0:0];
  _RAND_2376 = {1{`RANDOM}};
  _T_1826 = _RAND_2376[0:0];
  _RAND_2377 = {1{`RANDOM}};
  _T_1827 = _RAND_2377[0:0];
  _RAND_2378 = {1{`RANDOM}};
  _T_1828 = _RAND_2378[0:0];
  _RAND_2379 = {1{`RANDOM}};
  _T_1829 = _RAND_2379[0:0];
  _RAND_2380 = {1{`RANDOM}};
  _T_1830 = _RAND_2380[0:0];
  _RAND_2381 = {1{`RANDOM}};
  _T_1831 = _RAND_2381[0:0];
  _RAND_2382 = {1{`RANDOM}};
  _T_1832 = _RAND_2382[0:0];
  _RAND_2383 = {1{`RANDOM}};
  _T_1833 = _RAND_2383[0:0];
  _RAND_2384 = {1{`RANDOM}};
  _T_1834 = _RAND_2384[0:0];
  _RAND_2385 = {1{`RANDOM}};
  _T_1835 = _RAND_2385[0:0];
  _RAND_2386 = {1{`RANDOM}};
  _T_1836 = _RAND_2386[0:0];
  _RAND_2387 = {1{`RANDOM}};
  _T_1837 = _RAND_2387[0:0];
  _RAND_2388 = {1{`RANDOM}};
  _T_1838 = _RAND_2388[0:0];
  _RAND_2389 = {1{`RANDOM}};
  _T_1839 = _RAND_2389[0:0];
  _RAND_2390 = {1{`RANDOM}};
  _T_1840 = _RAND_2390[0:0];
  _RAND_2391 = {1{`RANDOM}};
  _T_1841 = _RAND_2391[0:0];
  _RAND_2392 = {1{`RANDOM}};
  _T_1842 = _RAND_2392[0:0];
  _RAND_2393 = {1{`RANDOM}};
  _T_1843 = _RAND_2393[0:0];
  _RAND_2394 = {1{`RANDOM}};
  _T_1844 = _RAND_2394[0:0];
  _RAND_2395 = {1{`RANDOM}};
  _T_1845 = _RAND_2395[0:0];
  _RAND_2396 = {1{`RANDOM}};
  _T_1846 = _RAND_2396[0:0];
  _RAND_2397 = {1{`RANDOM}};
  _T_1847 = _RAND_2397[0:0];
  _RAND_2398 = {1{`RANDOM}};
  _T_1848 = _RAND_2398[0:0];
  _RAND_2399 = {1{`RANDOM}};
  _T_1849 = _RAND_2399[0:0];
  _RAND_2400 = {1{`RANDOM}};
  _T_1850 = _RAND_2400[0:0];
  _RAND_2401 = {1{`RANDOM}};
  _T_1851 = _RAND_2401[0:0];
  _RAND_2402 = {1{`RANDOM}};
  _T_1852 = _RAND_2402[0:0];
  _RAND_2403 = {1{`RANDOM}};
  _T_1853 = _RAND_2403[0:0];
  _RAND_2404 = {1{`RANDOM}};
  _T_1854 = _RAND_2404[0:0];
  _RAND_2405 = {1{`RANDOM}};
  _T_1855 = _RAND_2405[0:0];
  _RAND_2406 = {1{`RANDOM}};
  _T_1856 = _RAND_2406[0:0];
  _RAND_2407 = {1{`RANDOM}};
  _T_1857 = _RAND_2407[0:0];
  _RAND_2408 = {1{`RANDOM}};
  _T_1858 = _RAND_2408[0:0];
  _RAND_2409 = {1{`RANDOM}};
  _T_1859 = _RAND_2409[0:0];
  _RAND_2410 = {1{`RANDOM}};
  _T_1860 = _RAND_2410[0:0];
  _RAND_2411 = {1{`RANDOM}};
  _T_1861 = _RAND_2411[0:0];
  _RAND_2412 = {1{`RANDOM}};
  _T_1862 = _RAND_2412[0:0];
  _RAND_2413 = {1{`RANDOM}};
  _T_1863 = _RAND_2413[0:0];
  _RAND_2414 = {1{`RANDOM}};
  _T_1864 = _RAND_2414[0:0];
  _RAND_2415 = {1{`RANDOM}};
  _T_1865 = _RAND_2415[0:0];
  _RAND_2416 = {1{`RANDOM}};
  _T_1866 = _RAND_2416[0:0];
  _RAND_2417 = {1{`RANDOM}};
  _T_1867 = _RAND_2417[0:0];
  _RAND_2418 = {1{`RANDOM}};
  _T_1868 = _RAND_2418[0:0];
  _RAND_2419 = {1{`RANDOM}};
  _T_1869 = _RAND_2419[0:0];
  _RAND_2420 = {1{`RANDOM}};
  _T_1870 = _RAND_2420[0:0];
  _RAND_2421 = {1{`RANDOM}};
  _T_1871 = _RAND_2421[0:0];
  _RAND_2422 = {1{`RANDOM}};
  _T_1872 = _RAND_2422[0:0];
  _RAND_2423 = {1{`RANDOM}};
  _T_1873 = _RAND_2423[0:0];
  _RAND_2424 = {1{`RANDOM}};
  _T_1874 = _RAND_2424[0:0];
  _RAND_2425 = {1{`RANDOM}};
  _T_1875 = _RAND_2425[0:0];
  _RAND_2426 = {1{`RANDOM}};
  _T_1876 = _RAND_2426[0:0];
  _RAND_2427 = {1{`RANDOM}};
  _T_1877 = _RAND_2427[0:0];
  _RAND_2428 = {1{`RANDOM}};
  _T_1878 = _RAND_2428[0:0];
  _RAND_2429 = {1{`RANDOM}};
  _T_1879 = _RAND_2429[0:0];
  _RAND_2430 = {1{`RANDOM}};
  _T_1880 = _RAND_2430[0:0];
  _RAND_2431 = {1{`RANDOM}};
  _T_1881 = _RAND_2431[0:0];
  _RAND_2432 = {1{`RANDOM}};
  _T_1882 = _RAND_2432[0:0];
  _RAND_2433 = {1{`RANDOM}};
  _T_1883 = _RAND_2433[0:0];
  _RAND_2434 = {1{`RANDOM}};
  _T_1884 = _RAND_2434[0:0];
  _RAND_2435 = {1{`RANDOM}};
  _T_1885 = _RAND_2435[0:0];
  _RAND_2436 = {1{`RANDOM}};
  _T_1886 = _RAND_2436[0:0];
  _RAND_2437 = {1{`RANDOM}};
  _T_1887 = _RAND_2437[0:0];
  _RAND_2438 = {1{`RANDOM}};
  _T_1888 = _RAND_2438[0:0];
  _RAND_2439 = {1{`RANDOM}};
  _T_1889 = _RAND_2439[0:0];
  _RAND_2440 = {1{`RANDOM}};
  _T_1890 = _RAND_2440[0:0];
  _RAND_2441 = {1{`RANDOM}};
  _T_1891 = _RAND_2441[0:0];
  _RAND_2442 = {1{`RANDOM}};
  _T_1892 = _RAND_2442[0:0];
  _RAND_2443 = {1{`RANDOM}};
  _T_1893 = _RAND_2443[0:0];
  _RAND_2444 = {1{`RANDOM}};
  _T_1894 = _RAND_2444[0:0];
  _RAND_2445 = {1{`RANDOM}};
  _T_1895 = _RAND_2445[0:0];
  _RAND_2446 = {1{`RANDOM}};
  _T_1896 = _RAND_2446[0:0];
  _RAND_2447 = {1{`RANDOM}};
  _T_1897 = _RAND_2447[0:0];
  _RAND_2448 = {1{`RANDOM}};
  _T_1898 = _RAND_2448[0:0];
  _RAND_2449 = {1{`RANDOM}};
  _T_1899 = _RAND_2449[0:0];
  _RAND_2450 = {1{`RANDOM}};
  _T_1900 = _RAND_2450[0:0];
  _RAND_2451 = {1{`RANDOM}};
  _T_1901 = _RAND_2451[0:0];
  _RAND_2452 = {1{`RANDOM}};
  _T_1902 = _RAND_2452[0:0];
  _RAND_2453 = {1{`RANDOM}};
  _T_1903 = _RAND_2453[0:0];
  _RAND_2454 = {1{`RANDOM}};
  _T_1904 = _RAND_2454[0:0];
  _RAND_2455 = {1{`RANDOM}};
  _T_1905 = _RAND_2455[0:0];
  _RAND_2456 = {1{`RANDOM}};
  _T_1906 = _RAND_2456[0:0];
  _RAND_2457 = {1{`RANDOM}};
  _T_1907 = _RAND_2457[0:0];
  _RAND_2458 = {1{`RANDOM}};
  _T_1908 = _RAND_2458[0:0];
  _RAND_2459 = {1{`RANDOM}};
  _T_1909 = _RAND_2459[0:0];
  _RAND_2460 = {1{`RANDOM}};
  _T_1910 = _RAND_2460[0:0];
  _RAND_2461 = {1{`RANDOM}};
  _T_1911 = _RAND_2461[0:0];
  _RAND_2462 = {1{`RANDOM}};
  _T_1912 = _RAND_2462[0:0];
  _RAND_2463 = {1{`RANDOM}};
  _T_1913 = _RAND_2463[0:0];
  _RAND_2464 = {1{`RANDOM}};
  _T_1914 = _RAND_2464[0:0];
  _RAND_2465 = {1{`RANDOM}};
  _T_1915 = _RAND_2465[0:0];
  _RAND_2466 = {1{`RANDOM}};
  _T_1916 = _RAND_2466[0:0];
  _RAND_2467 = {1{`RANDOM}};
  _T_1917 = _RAND_2467[0:0];
  _RAND_2468 = {1{`RANDOM}};
  _T_1918 = _RAND_2468[0:0];
  _RAND_2469 = {1{`RANDOM}};
  _T_1919 = _RAND_2469[0:0];
  _RAND_2470 = {1{`RANDOM}};
  _T_1920 = _RAND_2470[0:0];
  _RAND_2471 = {1{`RANDOM}};
  _T_1921 = _RAND_2471[0:0];
  _RAND_2472 = {1{`RANDOM}};
  _T_1922 = _RAND_2472[0:0];
  _RAND_2473 = {1{`RANDOM}};
  _T_1923 = _RAND_2473[0:0];
  _RAND_2474 = {1{`RANDOM}};
  _T_1924 = _RAND_2474[0:0];
  _RAND_2475 = {1{`RANDOM}};
  _T_1925 = _RAND_2475[0:0];
  _RAND_2476 = {1{`RANDOM}};
  _T_1926 = _RAND_2476[0:0];
  _RAND_2477 = {1{`RANDOM}};
  _T_1927 = _RAND_2477[0:0];
  _RAND_2478 = {1{`RANDOM}};
  _T_1928 = _RAND_2478[0:0];
  _RAND_2479 = {1{`RANDOM}};
  _T_1929 = _RAND_2479[0:0];
  _RAND_2480 = {1{`RANDOM}};
  _T_1930 = _RAND_2480[0:0];
  _RAND_2481 = {1{`RANDOM}};
  _T_1931 = _RAND_2481[0:0];
  _RAND_2482 = {1{`RANDOM}};
  _T_1932 = _RAND_2482[0:0];
  _RAND_2483 = {1{`RANDOM}};
  _T_1933 = _RAND_2483[0:0];
  _RAND_2484 = {1{`RANDOM}};
  _T_1934 = _RAND_2484[0:0];
  _RAND_2485 = {1{`RANDOM}};
  _T_1935 = _RAND_2485[0:0];
  _RAND_2486 = {1{`RANDOM}};
  _T_1936 = _RAND_2486[0:0];
  _RAND_2487 = {1{`RANDOM}};
  _T_1937 = _RAND_2487[0:0];
  _RAND_2488 = {1{`RANDOM}};
  _T_1938 = _RAND_2488[0:0];
  _RAND_2489 = {1{`RANDOM}};
  _T_1939 = _RAND_2489[0:0];
  _RAND_2490 = {1{`RANDOM}};
  _T_1940 = _RAND_2490[0:0];
  _RAND_2491 = {1{`RANDOM}};
  _T_1941 = _RAND_2491[0:0];
  _RAND_2492 = {1{`RANDOM}};
  _T_1942 = _RAND_2492[0:0];
  _RAND_2493 = {1{`RANDOM}};
  _T_1943 = _RAND_2493[0:0];
  _RAND_2494 = {1{`RANDOM}};
  _T_1944 = _RAND_2494[0:0];
  _RAND_2495 = {1{`RANDOM}};
  _T_1945 = _RAND_2495[0:0];
  _RAND_2496 = {1{`RANDOM}};
  _T_1946 = _RAND_2496[0:0];
  _RAND_2497 = {1{`RANDOM}};
  _T_1947 = _RAND_2497[0:0];
  _RAND_2498 = {1{`RANDOM}};
  _T_1948 = _RAND_2498[0:0];
  _RAND_2499 = {1{`RANDOM}};
  _T_1949 = _RAND_2499[0:0];
  _RAND_2500 = {1{`RANDOM}};
  _T_1950 = _RAND_2500[0:0];
  _RAND_2501 = {1{`RANDOM}};
  _T_1951 = _RAND_2501[0:0];
  _RAND_2502 = {1{`RANDOM}};
  _T_1952 = _RAND_2502[0:0];
  _RAND_2503 = {1{`RANDOM}};
  _T_1953 = _RAND_2503[0:0];
  _RAND_2504 = {1{`RANDOM}};
  _T_1954 = _RAND_2504[0:0];
  _RAND_2505 = {1{`RANDOM}};
  _T_1955 = _RAND_2505[0:0];
  _RAND_2506 = {1{`RANDOM}};
  _T_1956 = _RAND_2506[0:0];
  _RAND_2507 = {1{`RANDOM}};
  _T_1957 = _RAND_2507[0:0];
  _RAND_2508 = {1{`RANDOM}};
  _T_1958 = _RAND_2508[0:0];
  _RAND_2509 = {1{`RANDOM}};
  _T_1959 = _RAND_2509[0:0];
  _RAND_2510 = {1{`RANDOM}};
  _T_1960 = _RAND_2510[0:0];
  _RAND_2511 = {1{`RANDOM}};
  _T_1961 = _RAND_2511[0:0];
  _RAND_2512 = {1{`RANDOM}};
  _T_1962 = _RAND_2512[0:0];
  _RAND_2513 = {1{`RANDOM}};
  _T_1963 = _RAND_2513[0:0];
  _RAND_2514 = {1{`RANDOM}};
  _T_1964 = _RAND_2514[0:0];
  _RAND_2515 = {1{`RANDOM}};
  _T_1965 = _RAND_2515[0:0];
  _RAND_2516 = {1{`RANDOM}};
  _T_1966 = _RAND_2516[0:0];
  _RAND_2517 = {1{`RANDOM}};
  _T_1967 = _RAND_2517[0:0];
  _RAND_2518 = {1{`RANDOM}};
  _T_1968 = _RAND_2518[0:0];
  _RAND_2519 = {1{`RANDOM}};
  _T_1969 = _RAND_2519[0:0];
  _RAND_2520 = {1{`RANDOM}};
  _T_1970 = _RAND_2520[0:0];
  _RAND_2521 = {1{`RANDOM}};
  _T_1971 = _RAND_2521[0:0];
  _RAND_2522 = {1{`RANDOM}};
  _T_1972 = _RAND_2522[0:0];
  _RAND_2523 = {1{`RANDOM}};
  _T_1973 = _RAND_2523[0:0];
  _RAND_2524 = {1{`RANDOM}};
  _T_1974 = _RAND_2524[0:0];
  _RAND_2525 = {1{`RANDOM}};
  _T_1975 = _RAND_2525[0:0];
  _RAND_2526 = {1{`RANDOM}};
  _T_1976 = _RAND_2526[0:0];
  _RAND_2527 = {1{`RANDOM}};
  _T_1977 = _RAND_2527[0:0];
  _RAND_2528 = {1{`RANDOM}};
  _T_1978 = _RAND_2528[0:0];
  _RAND_2529 = {1{`RANDOM}};
  _T_1979 = _RAND_2529[0:0];
  _RAND_2530 = {1{`RANDOM}};
  _T_1980 = _RAND_2530[0:0];
  _RAND_2531 = {1{`RANDOM}};
  _T_1981 = _RAND_2531[0:0];
  _RAND_2532 = {1{`RANDOM}};
  _T_1982 = _RAND_2532[0:0];
  _RAND_2533 = {1{`RANDOM}};
  _T_1983 = _RAND_2533[0:0];
  _RAND_2534 = {1{`RANDOM}};
  _T_1984 = _RAND_2534[0:0];
  _RAND_2535 = {1{`RANDOM}};
  _T_1985 = _RAND_2535[0:0];
  _RAND_2536 = {1{`RANDOM}};
  _T_1986 = _RAND_2536[0:0];
  _RAND_2537 = {1{`RANDOM}};
  _T_1987 = _RAND_2537[0:0];
  _RAND_2538 = {1{`RANDOM}};
  _T_1988 = _RAND_2538[0:0];
  _RAND_2539 = {1{`RANDOM}};
  _T_1989 = _RAND_2539[0:0];
  _RAND_2540 = {1{`RANDOM}};
  _T_1990 = _RAND_2540[0:0];
  _RAND_2541 = {1{`RANDOM}};
  _T_1991 = _RAND_2541[0:0];
  _RAND_2542 = {1{`RANDOM}};
  _T_1992 = _RAND_2542[0:0];
  _RAND_2543 = {1{`RANDOM}};
  _T_1993 = _RAND_2543[0:0];
  _RAND_2544 = {1{`RANDOM}};
  _T_1994 = _RAND_2544[0:0];
  _RAND_2545 = {1{`RANDOM}};
  _T_1995 = _RAND_2545[0:0];
  _RAND_2546 = {1{`RANDOM}};
  _T_1996 = _RAND_2546[0:0];
  _RAND_2547 = {1{`RANDOM}};
  _T_1997 = _RAND_2547[0:0];
  _RAND_2548 = {1{`RANDOM}};
  _T_1998 = _RAND_2548[0:0];
  _RAND_2549 = {1{`RANDOM}};
  _T_1999 = _RAND_2549[0:0];
  _RAND_2550 = {1{`RANDOM}};
  _T_2000 = _RAND_2550[0:0];
  _RAND_2551 = {1{`RANDOM}};
  _T_2001 = _RAND_2551[0:0];
  _RAND_2552 = {1{`RANDOM}};
  _T_2002 = _RAND_2552[0:0];
  _RAND_2553 = {1{`RANDOM}};
  _T_2003 = _RAND_2553[0:0];
  _RAND_2554 = {1{`RANDOM}};
  _T_2004 = _RAND_2554[0:0];
  _RAND_2555 = {1{`RANDOM}};
  _T_2005 = _RAND_2555[0:0];
  _RAND_2556 = {1{`RANDOM}};
  _T_2006 = _RAND_2556[0:0];
  _RAND_2557 = {1{`RANDOM}};
  _T_2007 = _RAND_2557[0:0];
  _RAND_2558 = {1{`RANDOM}};
  _T_2008 = _RAND_2558[0:0];
  _RAND_2559 = {1{`RANDOM}};
  _T_2009 = _RAND_2559[0:0];
  _RAND_2560 = {1{`RANDOM}};
  _T_2010 = _RAND_2560[0:0];
  _RAND_2561 = {1{`RANDOM}};
  _T_2011 = _RAND_2561[0:0];
  _RAND_2562 = {1{`RANDOM}};
  _T_2012 = _RAND_2562[0:0];
  _RAND_2563 = {1{`RANDOM}};
  _T_2013 = _RAND_2563[0:0];
  _RAND_2564 = {1{`RANDOM}};
  _T_2014 = _RAND_2564[0:0];
  _RAND_2565 = {1{`RANDOM}};
  _T_2015 = _RAND_2565[0:0];
  _RAND_2566 = {1{`RANDOM}};
  _T_2016 = _RAND_2566[0:0];
  _RAND_2567 = {1{`RANDOM}};
  _T_2017 = _RAND_2567[0:0];
  _RAND_2568 = {1{`RANDOM}};
  _T_2018 = _RAND_2568[0:0];
  _RAND_2569 = {1{`RANDOM}};
  _T_2019 = _RAND_2569[0:0];
  _RAND_2570 = {1{`RANDOM}};
  _T_2020 = _RAND_2570[0:0];
  _RAND_2571 = {1{`RANDOM}};
  _T_2021 = _RAND_2571[0:0];
  _RAND_2572 = {1{`RANDOM}};
  _T_2022 = _RAND_2572[0:0];
  _RAND_2573 = {1{`RANDOM}};
  _T_2023 = _RAND_2573[0:0];
  _RAND_2574 = {1{`RANDOM}};
  _T_2024 = _RAND_2574[0:0];
  _RAND_2575 = {1{`RANDOM}};
  _T_2025 = _RAND_2575[0:0];
  _RAND_2576 = {1{`RANDOM}};
  _T_2026 = _RAND_2576[0:0];
  _RAND_2577 = {1{`RANDOM}};
  _T_2027 = _RAND_2577[0:0];
  _RAND_2578 = {1{`RANDOM}};
  _T_2028 = _RAND_2578[0:0];
  _RAND_2579 = {1{`RANDOM}};
  _T_2029 = _RAND_2579[0:0];
  _RAND_2580 = {1{`RANDOM}};
  _T_2030 = _RAND_2580[0:0];
  _RAND_2581 = {1{`RANDOM}};
  _T_2031 = _RAND_2581[0:0];
  _RAND_2582 = {1{`RANDOM}};
  _T_2032 = _RAND_2582[0:0];
  _RAND_2583 = {1{`RANDOM}};
  _T_2033 = _RAND_2583[0:0];
  _RAND_2584 = {1{`RANDOM}};
  _T_2034 = _RAND_2584[0:0];
  _RAND_2585 = {1{`RANDOM}};
  _T_2035 = _RAND_2585[0:0];
  _RAND_2586 = {1{`RANDOM}};
  _T_2036 = _RAND_2586[0:0];
  _RAND_2587 = {1{`RANDOM}};
  _T_2037 = _RAND_2587[0:0];
  _RAND_2588 = {1{`RANDOM}};
  _T_2038 = _RAND_2588[0:0];
  _RAND_2589 = {1{`RANDOM}};
  _T_2039 = _RAND_2589[0:0];
  _RAND_2590 = {1{`RANDOM}};
  _T_2040 = _RAND_2590[0:0];
  _RAND_2591 = {1{`RANDOM}};
  _T_2041 = _RAND_2591[0:0];
  _RAND_2592 = {1{`RANDOM}};
  _T_2042 = _RAND_2592[0:0];
  _RAND_2593 = {1{`RANDOM}};
  _T_2043 = _RAND_2593[0:0];
  _RAND_2594 = {1{`RANDOM}};
  _T_2044 = _RAND_2594[0:0];
  _RAND_2595 = {1{`RANDOM}};
  _T_2045 = _RAND_2595[0:0];
  _RAND_2596 = {1{`RANDOM}};
  _T_2046 = _RAND_2596[0:0];
  _RAND_2597 = {1{`RANDOM}};
  _T_2047 = _RAND_2597[0:0];
  _RAND_2598 = {1{`RANDOM}};
  _T_2048 = _RAND_2598[0:0];
  _RAND_2599 = {1{`RANDOM}};
  _T_2049 = _RAND_2599[0:0];
  _RAND_2600 = {1{`RANDOM}};
  _T_2050 = _RAND_2600[0:0];
  _RAND_2601 = {1{`RANDOM}};
  _T_2051 = _RAND_2601[0:0];
  _RAND_2602 = {1{`RANDOM}};
  _T_2052 = _RAND_2602[0:0];
  _RAND_2603 = {1{`RANDOM}};
  _T_2053 = _RAND_2603[0:0];
  _RAND_2604 = {1{`RANDOM}};
  _T_2054 = _RAND_2604[0:0];
  _RAND_2605 = {1{`RANDOM}};
  _T_2055 = _RAND_2605[0:0];
  _RAND_2606 = {1{`RANDOM}};
  _T_2056 = _RAND_2606[0:0];
  _RAND_2607 = {1{`RANDOM}};
  _T_2057 = _RAND_2607[0:0];
  _RAND_2608 = {1{`RANDOM}};
  _T_2058 = _RAND_2608[0:0];
  _RAND_2609 = {1{`RANDOM}};
  _T_2059 = _RAND_2609[0:0];
  _RAND_2610 = {1{`RANDOM}};
  _T_2060 = _RAND_2610[0:0];
  _RAND_2611 = {1{`RANDOM}};
  _T_2061 = _RAND_2611[0:0];
  _RAND_2612 = {1{`RANDOM}};
  _T_2062 = _RAND_2612[0:0];
  _RAND_2613 = {1{`RANDOM}};
  _T_2063 = _RAND_2613[0:0];
  _RAND_2614 = {1{`RANDOM}};
  _T_2064 = _RAND_2614[0:0];
  _RAND_2615 = {1{`RANDOM}};
  _T_2065 = _RAND_2615[0:0];
  _RAND_2616 = {1{`RANDOM}};
  _T_2066 = _RAND_2616[0:0];
  _RAND_2617 = {1{`RANDOM}};
  _T_2067 = _RAND_2617[0:0];
  _RAND_2618 = {1{`RANDOM}};
  _T_2068 = _RAND_2618[0:0];
  _RAND_2619 = {1{`RANDOM}};
  _T_2069 = _RAND_2619[0:0];
  _RAND_2620 = {1{`RANDOM}};
  _T_2070 = _RAND_2620[0:0];
  _RAND_2621 = {1{`RANDOM}};
  _T_2071 = _RAND_2621[0:0];
  _RAND_2622 = {1{`RANDOM}};
  _T_2072 = _RAND_2622[0:0];
  _RAND_2623 = {1{`RANDOM}};
  _T_2073 = _RAND_2623[0:0];
  _RAND_2624 = {1{`RANDOM}};
  _T_2074 = _RAND_2624[0:0];
  _RAND_2625 = {1{`RANDOM}};
  _T_2075 = _RAND_2625[0:0];
  _RAND_2626 = {1{`RANDOM}};
  _T_2076 = _RAND_2626[0:0];
  _RAND_2627 = {1{`RANDOM}};
  _T_2077 = _RAND_2627[0:0];
  _RAND_2628 = {1{`RANDOM}};
  _T_2078 = _RAND_2628[0:0];
  _RAND_2629 = {1{`RANDOM}};
  _T_2079 = _RAND_2629[0:0];
  _RAND_2630 = {1{`RANDOM}};
  _T_2080 = _RAND_2630[0:0];
  _RAND_2631 = {1{`RANDOM}};
  _T_2081 = _RAND_2631[0:0];
  _RAND_2632 = {1{`RANDOM}};
  _T_2082 = _RAND_2632[0:0];
  _RAND_2633 = {1{`RANDOM}};
  _T_2083 = _RAND_2633[0:0];
  _RAND_2634 = {1{`RANDOM}};
  _T_2084 = _RAND_2634[0:0];
  _RAND_2635 = {1{`RANDOM}};
  _T_2085 = _RAND_2635[0:0];
  _RAND_2636 = {1{`RANDOM}};
  _T_2086 = _RAND_2636[0:0];
  _RAND_2637 = {1{`RANDOM}};
  _T_2087 = _RAND_2637[0:0];
  _RAND_2638 = {1{`RANDOM}};
  _T_2088 = _RAND_2638[0:0];
  _RAND_2639 = {1{`RANDOM}};
  _T_2089 = _RAND_2639[0:0];
  _RAND_2640 = {1{`RANDOM}};
  _T_2090 = _RAND_2640[0:0];
  _RAND_2641 = {1{`RANDOM}};
  _T_2091 = _RAND_2641[0:0];
  _RAND_2642 = {1{`RANDOM}};
  _T_2092 = _RAND_2642[0:0];
  _RAND_2643 = {1{`RANDOM}};
  _T_2093 = _RAND_2643[0:0];
  _RAND_2644 = {1{`RANDOM}};
  _T_2094 = _RAND_2644[0:0];
  _RAND_2645 = {1{`RANDOM}};
  _T_2095 = _RAND_2645[0:0];
  _RAND_2646 = {1{`RANDOM}};
  _T_2096 = _RAND_2646[0:0];
  _RAND_2647 = {1{`RANDOM}};
  _T_2097 = _RAND_2647[0:0];
  _RAND_2648 = {1{`RANDOM}};
  _T_2098 = _RAND_2648[0:0];
  _RAND_2649 = {1{`RANDOM}};
  _T_2099 = _RAND_2649[0:0];
  _RAND_2650 = {1{`RANDOM}};
  _T_2100 = _RAND_2650[0:0];
  _RAND_2651 = {1{`RANDOM}};
  _T_2101 = _RAND_2651[0:0];
  _RAND_2652 = {1{`RANDOM}};
  _T_2102 = _RAND_2652[0:0];
  _RAND_2653 = {1{`RANDOM}};
  _T_2103 = _RAND_2653[0:0];
  _RAND_2654 = {1{`RANDOM}};
  _T_2104 = _RAND_2654[0:0];
  _RAND_2655 = {1{`RANDOM}};
  _T_2105 = _RAND_2655[0:0];
  _RAND_2656 = {1{`RANDOM}};
  _T_2106 = _RAND_2656[0:0];
  _RAND_2657 = {1{`RANDOM}};
  _T_2107 = _RAND_2657[0:0];
  _RAND_2658 = {1{`RANDOM}};
  _T_2108 = _RAND_2658[0:0];
  _RAND_2659 = {1{`RANDOM}};
  _T_2109 = _RAND_2659[0:0];
  _RAND_2660 = {1{`RANDOM}};
  _T_2110 = _RAND_2660[0:0];
  _RAND_2661 = {1{`RANDOM}};
  _T_2111 = _RAND_2661[0:0];
  _RAND_2662 = {1{`RANDOM}};
  _T_2112 = _RAND_2662[0:0];
  _RAND_2663 = {1{`RANDOM}};
  _T_2113 = _RAND_2663[0:0];
  _RAND_2664 = {1{`RANDOM}};
  _T_2114 = _RAND_2664[0:0];
  _RAND_2665 = {1{`RANDOM}};
  _T_2115 = _RAND_2665[0:0];
  _RAND_2666 = {1{`RANDOM}};
  _T_2116 = _RAND_2666[0:0];
  _RAND_2667 = {1{`RANDOM}};
  _T_2117 = _RAND_2667[0:0];
  _RAND_2668 = {1{`RANDOM}};
  _T_2118 = _RAND_2668[0:0];
  _RAND_2669 = {1{`RANDOM}};
  _T_2119 = _RAND_2669[0:0];
  _RAND_2670 = {1{`RANDOM}};
  _T_2120 = _RAND_2670[0:0];
  _RAND_2671 = {1{`RANDOM}};
  _T_2121 = _RAND_2671[0:0];
  _RAND_2672 = {1{`RANDOM}};
  _T_2122 = _RAND_2672[0:0];
  _RAND_2673 = {1{`RANDOM}};
  _T_2123 = _RAND_2673[0:0];
  _RAND_2674 = {1{`RANDOM}};
  _T_2124 = _RAND_2674[0:0];
  _RAND_2675 = {1{`RANDOM}};
  _T_2125 = _RAND_2675[0:0];
  _RAND_2676 = {1{`RANDOM}};
  _T_2126 = _RAND_2676[0:0];
  _RAND_2677 = {1{`RANDOM}};
  _T_2127 = _RAND_2677[0:0];
  _RAND_2678 = {1{`RANDOM}};
  _T_2128 = _RAND_2678[0:0];
  _RAND_2679 = {1{`RANDOM}};
  _T_2129 = _RAND_2679[0:0];
  _RAND_2680 = {1{`RANDOM}};
  _T_2130 = _RAND_2680[0:0];
  _RAND_2681 = {1{`RANDOM}};
  _T_2131 = _RAND_2681[0:0];
  _RAND_2682 = {1{`RANDOM}};
  _T_2132 = _RAND_2682[0:0];
  _RAND_2683 = {1{`RANDOM}};
  _T_2133 = _RAND_2683[0:0];
  _RAND_2684 = {1{`RANDOM}};
  _T_2134 = _RAND_2684[0:0];
  _RAND_2685 = {1{`RANDOM}};
  _T_2135 = _RAND_2685[0:0];
  _RAND_2686 = {1{`RANDOM}};
  _T_2136 = _RAND_2686[0:0];
  _RAND_2687 = {1{`RANDOM}};
  _T_2137 = _RAND_2687[0:0];
  _RAND_2688 = {1{`RANDOM}};
  _T_2138 = _RAND_2688[0:0];
  _RAND_2689 = {1{`RANDOM}};
  _T_2139 = _RAND_2689[0:0];
  _RAND_2690 = {1{`RANDOM}};
  _T_2140 = _RAND_2690[0:0];
  _RAND_2691 = {1{`RANDOM}};
  _T_2141 = _RAND_2691[0:0];
  _RAND_2692 = {1{`RANDOM}};
  _T_2142 = _RAND_2692[0:0];
  _RAND_2693 = {1{`RANDOM}};
  _T_2143 = _RAND_2693[0:0];
  _RAND_2694 = {1{`RANDOM}};
  _T_2144 = _RAND_2694[0:0];
  _RAND_2695 = {1{`RANDOM}};
  _T_2145 = _RAND_2695[0:0];
  _RAND_2696 = {1{`RANDOM}};
  _T_2146 = _RAND_2696[0:0];
  _RAND_2697 = {1{`RANDOM}};
  _T_2147 = _RAND_2697[0:0];
  _RAND_2698 = {1{`RANDOM}};
  _T_2148 = _RAND_2698[0:0];
  _RAND_2699 = {1{`RANDOM}};
  _T_2149 = _RAND_2699[0:0];
  _RAND_2700 = {1{`RANDOM}};
  _T_2150 = _RAND_2700[0:0];
  _RAND_2701 = {1{`RANDOM}};
  _T_2151 = _RAND_2701[0:0];
  _RAND_2702 = {1{`RANDOM}};
  _T_2152 = _RAND_2702[0:0];
  _RAND_2703 = {1{`RANDOM}};
  _T_2153 = _RAND_2703[0:0];
  _RAND_2704 = {1{`RANDOM}};
  _T_2154 = _RAND_2704[0:0];
  _RAND_2705 = {1{`RANDOM}};
  _T_2155 = _RAND_2705[0:0];
  _RAND_2706 = {1{`RANDOM}};
  _T_2156 = _RAND_2706[0:0];
  _RAND_2707 = {1{`RANDOM}};
  _T_2157 = _RAND_2707[0:0];
  _RAND_2708 = {1{`RANDOM}};
  _T_2158 = _RAND_2708[0:0];
  _RAND_2709 = {1{`RANDOM}};
  _T_2159 = _RAND_2709[0:0];
  _RAND_2710 = {1{`RANDOM}};
  _T_2160 = _RAND_2710[0:0];
  _RAND_2711 = {1{`RANDOM}};
  _T_2161 = _RAND_2711[0:0];
  _RAND_2712 = {1{`RANDOM}};
  _T_2162 = _RAND_2712[0:0];
  _RAND_2713 = {1{`RANDOM}};
  _T_2163 = _RAND_2713[0:0];
  _RAND_2714 = {1{`RANDOM}};
  _T_2164 = _RAND_2714[0:0];
  _RAND_2715 = {1{`RANDOM}};
  _T_2165 = _RAND_2715[0:0];
  _RAND_2716 = {1{`RANDOM}};
  _T_2166 = _RAND_2716[0:0];
  _RAND_2717 = {1{`RANDOM}};
  _T_2167 = _RAND_2717[0:0];
  _RAND_2718 = {1{`RANDOM}};
  _T_2168 = _RAND_2718[0:0];
  _RAND_2719 = {1{`RANDOM}};
  _T_2169 = _RAND_2719[0:0];
  _RAND_2720 = {1{`RANDOM}};
  _T_2170 = _RAND_2720[0:0];
  _RAND_2721 = {1{`RANDOM}};
  _T_2171 = _RAND_2721[0:0];
  _RAND_2722 = {1{`RANDOM}};
  _T_2172 = _RAND_2722[0:0];
  _RAND_2723 = {1{`RANDOM}};
  _T_2173 = _RAND_2723[0:0];
  _RAND_2724 = {1{`RANDOM}};
  _T_2174 = _RAND_2724[0:0];
  _RAND_2725 = {1{`RANDOM}};
  _T_2175 = _RAND_2725[0:0];
  _RAND_2726 = {1{`RANDOM}};
  _T_2176 = _RAND_2726[0:0];
  _RAND_2727 = {1{`RANDOM}};
  _T_2177 = _RAND_2727[0:0];
  _RAND_2728 = {1{`RANDOM}};
  _T_2178 = _RAND_2728[0:0];
  _RAND_2729 = {1{`RANDOM}};
  _T_2179 = _RAND_2729[0:0];
  _RAND_2730 = {1{`RANDOM}};
  _T_2180 = _RAND_2730[0:0];
  _RAND_2731 = {1{`RANDOM}};
  _T_2181 = _RAND_2731[0:0];
  _RAND_2732 = {1{`RANDOM}};
  _T_2182 = _RAND_2732[0:0];
  _RAND_2733 = {1{`RANDOM}};
  _T_2183 = _RAND_2733[0:0];
  _RAND_2734 = {1{`RANDOM}};
  _T_2184 = _RAND_2734[0:0];
  _RAND_2735 = {1{`RANDOM}};
  _T_2185 = _RAND_2735[0:0];
  _RAND_2736 = {1{`RANDOM}};
  _T_2186 = _RAND_2736[0:0];
  _RAND_2737 = {1{`RANDOM}};
  _T_2187 = _RAND_2737[0:0];
  _RAND_2738 = {1{`RANDOM}};
  _T_2188 = _RAND_2738[0:0];
  _RAND_2739 = {1{`RANDOM}};
  _T_2189 = _RAND_2739[0:0];
  _RAND_2740 = {1{`RANDOM}};
  _T_2190 = _RAND_2740[0:0];
  _RAND_2741 = {1{`RANDOM}};
  _T_2191 = _RAND_2741[0:0];
  _RAND_2742 = {1{`RANDOM}};
  _T_2192 = _RAND_2742[0:0];
  _RAND_2743 = {1{`RANDOM}};
  _T_2193 = _RAND_2743[0:0];
  _RAND_2744 = {1{`RANDOM}};
  _T_2194 = _RAND_2744[0:0];
  _RAND_2745 = {1{`RANDOM}};
  _T_2195 = _RAND_2745[0:0];
  _RAND_2746 = {1{`RANDOM}};
  _T_2196 = _RAND_2746[0:0];
  _RAND_2747 = {1{`RANDOM}};
  _T_2197 = _RAND_2747[0:0];
  _RAND_2748 = {1{`RANDOM}};
  _T_2198 = _RAND_2748[0:0];
  _RAND_2749 = {1{`RANDOM}};
  _T_2199 = _RAND_2749[0:0];
  _RAND_2750 = {1{`RANDOM}};
  _T_2200 = _RAND_2750[0:0];
  _RAND_2751 = {1{`RANDOM}};
  _T_2201 = _RAND_2751[0:0];
  _RAND_2752 = {1{`RANDOM}};
  _T_2202 = _RAND_2752[0:0];
  _RAND_2753 = {1{`RANDOM}};
  _T_2203 = _RAND_2753[0:0];
  _RAND_2754 = {1{`RANDOM}};
  _T_2204 = _RAND_2754[0:0];
  _RAND_2755 = {1{`RANDOM}};
  _T_2205 = _RAND_2755[0:0];
  _RAND_2756 = {1{`RANDOM}};
  _T_2206 = _RAND_2756[0:0];
  _RAND_2757 = {1{`RANDOM}};
  _T_2207 = _RAND_2757[0:0];
  _RAND_2758 = {1{`RANDOM}};
  _T_2208 = _RAND_2758[0:0];
  _RAND_2759 = {1{`RANDOM}};
  _T_2209 = _RAND_2759[0:0];
  _RAND_2760 = {1{`RANDOM}};
  _T_2210 = _RAND_2760[0:0];
  _RAND_2761 = {1{`RANDOM}};
  _T_2211 = _RAND_2761[0:0];
  _RAND_2762 = {1{`RANDOM}};
  _T_2212 = _RAND_2762[0:0];
  _RAND_2763 = {1{`RANDOM}};
  _T_2213 = _RAND_2763[0:0];
  _RAND_2764 = {1{`RANDOM}};
  _T_2214 = _RAND_2764[0:0];
  _RAND_2765 = {1{`RANDOM}};
  _T_2215 = _RAND_2765[0:0];
  _RAND_2766 = {1{`RANDOM}};
  _T_2216 = _RAND_2766[0:0];
  _RAND_2767 = {1{`RANDOM}};
  _T_2217 = _RAND_2767[0:0];
  _RAND_2768 = {1{`RANDOM}};
  _T_2218 = _RAND_2768[0:0];
  _RAND_2769 = {1{`RANDOM}};
  _T_2219 = _RAND_2769[0:0];
  _RAND_2770 = {1{`RANDOM}};
  _T_2220 = _RAND_2770[0:0];
  _RAND_2771 = {1{`RANDOM}};
  _T_2221 = _RAND_2771[0:0];
  _RAND_2772 = {1{`RANDOM}};
  _T_2222 = _RAND_2772[0:0];
  _RAND_2773 = {1{`RANDOM}};
  _T_2223 = _RAND_2773[0:0];
  _RAND_2774 = {1{`RANDOM}};
  _T_2224 = _RAND_2774[0:0];
  _RAND_2775 = {1{`RANDOM}};
  _T_2225 = _RAND_2775[0:0];
  _RAND_2776 = {1{`RANDOM}};
  _T_2226 = _RAND_2776[0:0];
  _RAND_2777 = {1{`RANDOM}};
  _T_2227 = _RAND_2777[0:0];
  _RAND_2778 = {1{`RANDOM}};
  _T_2228 = _RAND_2778[0:0];
  _RAND_2779 = {1{`RANDOM}};
  _T_2229 = _RAND_2779[0:0];
  _RAND_2780 = {1{`RANDOM}};
  _T_2230 = _RAND_2780[0:0];
  _RAND_2781 = {1{`RANDOM}};
  _T_2231 = _RAND_2781[0:0];
  _RAND_2782 = {1{`RANDOM}};
  _T_2232 = _RAND_2782[0:0];
  _RAND_2783 = {1{`RANDOM}};
  _T_2233 = _RAND_2783[0:0];
  _RAND_2784 = {1{`RANDOM}};
  _T_2234 = _RAND_2784[0:0];
  _RAND_2785 = {1{`RANDOM}};
  _T_2235 = _RAND_2785[0:0];
  _RAND_2786 = {1{`RANDOM}};
  _T_2236 = _RAND_2786[0:0];
  _RAND_2787 = {1{`RANDOM}};
  _T_2237 = _RAND_2787[0:0];
  _RAND_2788 = {1{`RANDOM}};
  _T_2238 = _RAND_2788[0:0];
  _RAND_2789 = {1{`RANDOM}};
  _T_2239 = _RAND_2789[0:0];
  _RAND_2790 = {1{`RANDOM}};
  _T_2240 = _RAND_2790[0:0];
  _RAND_2791 = {1{`RANDOM}};
  _T_2241 = _RAND_2791[0:0];
  _RAND_2792 = {1{`RANDOM}};
  _T_2242 = _RAND_2792[0:0];
  _RAND_2793 = {1{`RANDOM}};
  _T_2243 = _RAND_2793[0:0];
  _RAND_2794 = {1{`RANDOM}};
  _T_2244 = _RAND_2794[0:0];
  _RAND_2795 = {1{`RANDOM}};
  _T_2245 = _RAND_2795[0:0];
  _RAND_2796 = {1{`RANDOM}};
  _T_2246 = _RAND_2796[0:0];
  _RAND_2797 = {1{`RANDOM}};
  _T_2247 = _RAND_2797[0:0];
  _RAND_2798 = {1{`RANDOM}};
  _T_2248 = _RAND_2798[0:0];
  _RAND_2799 = {1{`RANDOM}};
  _T_2249 = _RAND_2799[0:0];
  _RAND_2800 = {1{`RANDOM}};
  _T_2250 = _RAND_2800[0:0];
  _RAND_2801 = {1{`RANDOM}};
  _T_2251 = _RAND_2801[0:0];
  _RAND_2802 = {1{`RANDOM}};
  _T_2252 = _RAND_2802[0:0];
  _RAND_2803 = {1{`RANDOM}};
  _T_2253 = _RAND_2803[0:0];
  _RAND_2804 = {1{`RANDOM}};
  _T_2254 = _RAND_2804[0:0];
  _RAND_2805 = {1{`RANDOM}};
  _T_2255 = _RAND_2805[0:0];
  _RAND_2806 = {1{`RANDOM}};
  _T_2256 = _RAND_2806[0:0];
  _RAND_2807 = {1{`RANDOM}};
  _T_2257 = _RAND_2807[0:0];
  _RAND_2808 = {1{`RANDOM}};
  _T_2258 = _RAND_2808[0:0];
  _RAND_2809 = {1{`RANDOM}};
  _T_2259 = _RAND_2809[0:0];
  _RAND_2810 = {1{`RANDOM}};
  _T_2260 = _RAND_2810[0:0];
  _RAND_2811 = {1{`RANDOM}};
  _T_2261 = _RAND_2811[0:0];
  _RAND_2812 = {1{`RANDOM}};
  _T_2262 = _RAND_2812[0:0];
  _RAND_2813 = {1{`RANDOM}};
  _T_2263 = _RAND_2813[0:0];
  _RAND_2814 = {1{`RANDOM}};
  _T_2264 = _RAND_2814[0:0];
  _RAND_2815 = {1{`RANDOM}};
  _T_2265 = _RAND_2815[0:0];
  _RAND_2816 = {1{`RANDOM}};
  _T_2266 = _RAND_2816[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 9'h0;
    end else if (io_din_valid) begin
      cnt <= _T_1;
    end
    _T_150_re <= io_dIn_re;
    _T_150_im <= io_dIn_im;
    _T_151_re <= _T_150_re;
    _T_151_im <= _T_150_im;
    _T_152_re <= _T_151_re;
    _T_152_im <= _T_151_im;
    _T_153_re <= _T_152_re;
    _T_153_im <= _T_152_im;
    _T_154_re <= _T_153_re;
    _T_154_im <= _T_153_im;
    _T_155_re <= _T_154_re;
    _T_155_im <= _T_154_im;
    _T_156_re <= _T_155_re;
    _T_156_im <= _T_155_im;
    _T_157_re <= _T_156_re;
    _T_157_im <= _T_156_im;
    _T_158_re <= _T_157_re;
    _T_158_im <= _T_157_im;
    _T_159_re <= _T_158_re;
    _T_159_im <= _T_158_im;
    _T_160_re <= _T_159_re;
    _T_160_im <= _T_159_im;
    _T_161_re <= _T_160_re;
    _T_161_im <= _T_160_im;
    _T_162_re <= _T_161_re;
    _T_162_im <= _T_161_im;
    _T_163_re <= _T_162_re;
    _T_163_im <= _T_162_im;
    _T_164_re <= _T_163_re;
    _T_164_im <= _T_163_im;
    _T_165_re <= _T_164_re;
    _T_165_im <= _T_164_im;
    _T_166_re <= _T_165_re;
    _T_166_im <= _T_165_im;
    _T_167_re <= _T_166_re;
    _T_167_im <= _T_166_im;
    _T_168_re <= _T_167_re;
    _T_168_im <= _T_167_im;
    _T_169_re <= _T_168_re;
    _T_169_im <= _T_168_im;
    _T_170_re <= _T_169_re;
    _T_170_im <= _T_169_im;
    _T_171_re <= _T_170_re;
    _T_171_im <= _T_170_im;
    _T_172_re <= _T_171_re;
    _T_172_im <= _T_171_im;
    _T_173_re <= _T_172_re;
    _T_173_im <= _T_172_im;
    _T_174_re <= _T_173_re;
    _T_174_im <= _T_173_im;
    _T_175_re <= _T_174_re;
    _T_175_im <= _T_174_im;
    _T_176_re <= _T_175_re;
    _T_176_im <= _T_175_im;
    _T_177_re <= _T_176_re;
    _T_177_im <= _T_176_im;
    _T_178_re <= _T_177_re;
    _T_178_im <= _T_177_im;
    _T_179_re <= _T_178_re;
    _T_179_im <= _T_178_im;
    _T_180_re <= _T_179_re;
    _T_180_im <= _T_179_im;
    _T_181_re <= _T_180_re;
    _T_181_im <= _T_180_im;
    _T_182_re <= _T_181_re;
    _T_182_im <= _T_181_im;
    _T_183_re <= _T_182_re;
    _T_183_im <= _T_182_im;
    _T_184_re <= _T_183_re;
    _T_184_im <= _T_183_im;
    _T_185_re <= _T_184_re;
    _T_185_im <= _T_184_im;
    _T_186_re <= _T_185_re;
    _T_186_im <= _T_185_im;
    _T_187_re <= _T_186_re;
    _T_187_im <= _T_186_im;
    _T_188_re <= _T_187_re;
    _T_188_im <= _T_187_im;
    _T_189_re <= _T_188_re;
    _T_189_im <= _T_188_im;
    _T_190_re <= _T_189_re;
    _T_190_im <= _T_189_im;
    _T_191_re <= _T_190_re;
    _T_191_im <= _T_190_im;
    _T_192_re <= _T_191_re;
    _T_192_im <= _T_191_im;
    _T_193_re <= _T_192_re;
    _T_193_im <= _T_192_im;
    _T_194_re <= _T_193_re;
    _T_194_im <= _T_193_im;
    _T_195_re <= _T_194_re;
    _T_195_im <= _T_194_im;
    _T_196_re <= _T_195_re;
    _T_196_im <= _T_195_im;
    _T_197_re <= _T_196_re;
    _T_197_im <= _T_196_im;
    _T_198_re <= _T_197_re;
    _T_198_im <= _T_197_im;
    _T_199_re <= _T_198_re;
    _T_199_im <= _T_198_im;
    _T_200_re <= _T_199_re;
    _T_200_im <= _T_199_im;
    _T_201_re <= _T_200_re;
    _T_201_im <= _T_200_im;
    _T_202_re <= _T_201_re;
    _T_202_im <= _T_201_im;
    _T_203_re <= _T_202_re;
    _T_203_im <= _T_202_im;
    _T_204_re <= _T_203_re;
    _T_204_im <= _T_203_im;
    _T_205_re <= _T_204_re;
    _T_205_im <= _T_204_im;
    _T_206_re <= _T_205_re;
    _T_206_im <= _T_205_im;
    _T_207_re <= _T_206_re;
    _T_207_im <= _T_206_im;
    _T_208_re <= _T_207_re;
    _T_208_im <= _T_207_im;
    _T_209_re <= _T_208_re;
    _T_209_im <= _T_208_im;
    _T_210_re <= _T_209_re;
    _T_210_im <= _T_209_im;
    _T_211_re <= _T_210_re;
    _T_211_im <= _T_210_im;
    _T_212_re <= _T_211_re;
    _T_212_im <= _T_211_im;
    _T_213_re <= _T_212_re;
    _T_213_im <= _T_212_im;
    _T_214_re <= _T_213_re;
    _T_214_im <= _T_213_im;
    _T_215_re <= _T_214_re;
    _T_215_im <= _T_214_im;
    _T_216_re <= _T_215_re;
    _T_216_im <= _T_215_im;
    _T_217_re <= _T_216_re;
    _T_217_im <= _T_216_im;
    _T_218_re <= _T_217_re;
    _T_218_im <= _T_217_im;
    _T_219_re <= _T_218_re;
    _T_219_im <= _T_218_im;
    _T_220_re <= _T_219_re;
    _T_220_im <= _T_219_im;
    _T_221_re <= _T_220_re;
    _T_221_im <= _T_220_im;
    _T_222_re <= _T_221_re;
    _T_222_im <= _T_221_im;
    _T_223_re <= _T_222_re;
    _T_223_im <= _T_222_im;
    _T_224_re <= _T_223_re;
    _T_224_im <= _T_223_im;
    _T_225_re <= _T_224_re;
    _T_225_im <= _T_224_im;
    _T_226_re <= _T_225_re;
    _T_226_im <= _T_225_im;
    _T_227_re <= _T_226_re;
    _T_227_im <= _T_226_im;
    _T_228_re <= _T_227_re;
    _T_228_im <= _T_227_im;
    _T_229_re <= _T_228_re;
    _T_229_im <= _T_228_im;
    _T_230_re <= _T_229_re;
    _T_230_im <= _T_229_im;
    _T_231_re <= _T_230_re;
    _T_231_im <= _T_230_im;
    _T_232_re <= _T_231_re;
    _T_232_im <= _T_231_im;
    _T_233_re <= _T_232_re;
    _T_233_im <= _T_232_im;
    _T_234_re <= _T_233_re;
    _T_234_im <= _T_233_im;
    _T_235_re <= _T_234_re;
    _T_235_im <= _T_234_im;
    _T_236_re <= _T_235_re;
    _T_236_im <= _T_235_im;
    _T_237_re <= _T_236_re;
    _T_237_im <= _T_236_im;
    _T_238_re <= _T_237_re;
    _T_238_im <= _T_237_im;
    _T_239_re <= _T_238_re;
    _T_239_im <= _T_238_im;
    _T_240_re <= _T_239_re;
    _T_240_im <= _T_239_im;
    _T_241_re <= _T_240_re;
    _T_241_im <= _T_240_im;
    _T_242_re <= _T_241_re;
    _T_242_im <= _T_241_im;
    _T_243_re <= _T_242_re;
    _T_243_im <= _T_242_im;
    _T_244_re <= _T_243_re;
    _T_244_im <= _T_243_im;
    _T_245_re <= _T_244_re;
    _T_245_im <= _T_244_im;
    _T_246_re <= _T_245_re;
    _T_246_im <= _T_245_im;
    _T_247_re <= _T_246_re;
    _T_247_im <= _T_246_im;
    _T_248_re <= _T_247_re;
    _T_248_im <= _T_247_im;
    _T_249_re <= _T_248_re;
    _T_249_im <= _T_248_im;
    _T_250_re <= _T_249_re;
    _T_250_im <= _T_249_im;
    _T_251_re <= _T_250_re;
    _T_251_im <= _T_250_im;
    _T_252_re <= _T_251_re;
    _T_252_im <= _T_251_im;
    _T_253_re <= _T_252_re;
    _T_253_im <= _T_252_im;
    _T_254_re <= _T_253_re;
    _T_254_im <= _T_253_im;
    _T_255_re <= _T_254_re;
    _T_255_im <= _T_254_im;
    _T_256_re <= _T_255_re;
    _T_256_im <= _T_255_im;
    _T_257_re <= _T_256_re;
    _T_257_im <= _T_256_im;
    _T_258_re <= _T_257_re;
    _T_258_im <= _T_257_im;
    _T_259_re <= _T_258_re;
    _T_259_im <= _T_258_im;
    _T_260_re <= _T_259_re;
    _T_260_im <= _T_259_im;
    _T_261_re <= _T_260_re;
    _T_261_im <= _T_260_im;
    _T_262_re <= _T_261_re;
    _T_262_im <= _T_261_im;
    _T_263_re <= _T_262_re;
    _T_263_im <= _T_262_im;
    _T_264_re <= _T_263_re;
    _T_264_im <= _T_263_im;
    _T_265_re <= _T_264_re;
    _T_265_im <= _T_264_im;
    _T_266_re <= _T_265_re;
    _T_266_im <= _T_265_im;
    _T_267_re <= _T_266_re;
    _T_267_im <= _T_266_im;
    _T_268_re <= _T_267_re;
    _T_268_im <= _T_267_im;
    _T_269_re <= _T_268_re;
    _T_269_im <= _T_268_im;
    _T_270_re <= _T_269_re;
    _T_270_im <= _T_269_im;
    _T_271_re <= _T_270_re;
    _T_271_im <= _T_270_im;
    _T_272_re <= _T_271_re;
    _T_272_im <= _T_271_im;
    _T_273_re <= _T_272_re;
    _T_273_im <= _T_272_im;
    _T_274_re <= _T_273_re;
    _T_274_im <= _T_273_im;
    _T_275_re <= _T_274_re;
    _T_275_im <= _T_274_im;
    _T_276_re <= _T_275_re;
    _T_276_im <= _T_275_im;
    _T_277_re <= _T_276_re;
    _T_277_im <= _T_276_im;
    _T_278_re <= _T_277_re;
    _T_278_im <= _T_277_im;
    _T_279_re <= _T_278_re;
    _T_279_im <= _T_278_im;
    _T_280_re <= _T_279_re;
    _T_280_im <= _T_279_im;
    _T_281_re <= _T_280_re;
    _T_281_im <= _T_280_im;
    _T_282_re <= _T_281_re;
    _T_282_im <= _T_281_im;
    _T_283_re <= _T_282_re;
    _T_283_im <= _T_282_im;
    _T_284_re <= _T_283_re;
    _T_284_im <= _T_283_im;
    _T_285_re <= _T_284_re;
    _T_285_im <= _T_284_im;
    _T_286_re <= _T_285_re;
    _T_286_im <= _T_285_im;
    _T_287_re <= _T_286_re;
    _T_287_im <= _T_286_im;
    _T_288_re <= _T_287_re;
    _T_288_im <= _T_287_im;
    _T_289_re <= _T_288_re;
    _T_289_im <= _T_288_im;
    _T_290_re <= _T_289_re;
    _T_290_im <= _T_289_im;
    _T_291_re <= _T_290_re;
    _T_291_im <= _T_290_im;
    _T_292_re <= _T_291_re;
    _T_292_im <= _T_291_im;
    _T_293_re <= _T_292_re;
    _T_293_im <= _T_292_im;
    _T_294_re <= _T_293_re;
    _T_294_im <= _T_293_im;
    _T_295_re <= _T_294_re;
    _T_295_im <= _T_294_im;
    _T_296_re <= _T_295_re;
    _T_296_im <= _T_295_im;
    _T_297_re <= _T_296_re;
    _T_297_im <= _T_296_im;
    _T_298_re <= _T_297_re;
    _T_298_im <= _T_297_im;
    _T_299_re <= _T_298_re;
    _T_299_im <= _T_298_im;
    _T_300_re <= _T_299_re;
    _T_300_im <= _T_299_im;
    _T_301_re <= _T_300_re;
    _T_301_im <= _T_300_im;
    _T_302_re <= _T_301_re;
    _T_302_im <= _T_301_im;
    _T_303_re <= _T_302_re;
    _T_303_im <= _T_302_im;
    _T_304_re <= _T_303_re;
    _T_304_im <= _T_303_im;
    _T_305_re <= _T_304_re;
    _T_305_im <= _T_304_im;
    _T_306_re <= _T_305_re;
    _T_306_im <= _T_305_im;
    _T_307_re <= _T_306_re;
    _T_307_im <= _T_306_im;
    _T_308_re <= _T_307_re;
    _T_308_im <= _T_307_im;
    _T_309_re <= _T_308_re;
    _T_309_im <= _T_308_im;
    _T_310_re <= _T_309_re;
    _T_310_im <= _T_309_im;
    _T_311_re <= _T_310_re;
    _T_311_im <= _T_310_im;
    _T_312_re <= _T_311_re;
    _T_312_im <= _T_311_im;
    _T_313_re <= _T_312_re;
    _T_313_im <= _T_312_im;
    _T_314_re <= _T_313_re;
    _T_314_im <= _T_313_im;
    _T_315_re <= _T_314_re;
    _T_315_im <= _T_314_im;
    _T_316_re <= _T_315_re;
    _T_316_im <= _T_315_im;
    _T_317_re <= _T_316_re;
    _T_317_im <= _T_316_im;
    _T_318_re <= _T_317_re;
    _T_318_im <= _T_317_im;
    _T_319_re <= _T_318_re;
    _T_319_im <= _T_318_im;
    _T_320_re <= _T_319_re;
    _T_320_im <= _T_319_im;
    _T_321_re <= _T_320_re;
    _T_321_im <= _T_320_im;
    _T_322_re <= _T_321_re;
    _T_322_im <= _T_321_im;
    _T_323_re <= _T_322_re;
    _T_323_im <= _T_322_im;
    _T_324_re <= _T_323_re;
    _T_324_im <= _T_323_im;
    _T_325_re <= _T_324_re;
    _T_325_im <= _T_324_im;
    _T_326_re <= _T_325_re;
    _T_326_im <= _T_325_im;
    _T_327_re <= _T_326_re;
    _T_327_im <= _T_326_im;
    _T_328_re <= _T_327_re;
    _T_328_im <= _T_327_im;
    _T_329_re <= _T_328_re;
    _T_329_im <= _T_328_im;
    _T_330_re <= _T_329_re;
    _T_330_im <= _T_329_im;
    _T_331_re <= _T_330_re;
    _T_331_im <= _T_330_im;
    _T_332_re <= _T_331_re;
    _T_332_im <= _T_331_im;
    _T_333_re <= _T_332_re;
    _T_333_im <= _T_332_im;
    _T_334_re <= _T_333_re;
    _T_334_im <= _T_333_im;
    _T_335_re <= _T_334_re;
    _T_335_im <= _T_334_im;
    _T_336_re <= _T_335_re;
    _T_336_im <= _T_335_im;
    _T_337_re <= _T_336_re;
    _T_337_im <= _T_336_im;
    _T_338_re <= _T_337_re;
    _T_338_im <= _T_337_im;
    _T_339_re <= _T_338_re;
    _T_339_im <= _T_338_im;
    _T_340_re <= _T_339_re;
    _T_340_im <= _T_339_im;
    _T_341_re <= _T_340_re;
    _T_341_im <= _T_340_im;
    _T_342_re <= _T_341_re;
    _T_342_im <= _T_341_im;
    _T_343_re <= _T_342_re;
    _T_343_im <= _T_342_im;
    _T_344_re <= _T_343_re;
    _T_344_im <= _T_343_im;
    _T_345_re <= _T_344_re;
    _T_345_im <= _T_344_im;
    _T_346_re <= _T_345_re;
    _T_346_im <= _T_345_im;
    _T_347_re <= _T_346_re;
    _T_347_im <= _T_346_im;
    _T_348_re <= _T_347_re;
    _T_348_im <= _T_347_im;
    _T_349_re <= _T_348_re;
    _T_349_im <= _T_348_im;
    _T_350_re <= _T_349_re;
    _T_350_im <= _T_349_im;
    _T_351_re <= _T_350_re;
    _T_351_im <= _T_350_im;
    _T_352_re <= _T_351_re;
    _T_352_im <= _T_351_im;
    _T_353_re <= _T_352_re;
    _T_353_im <= _T_352_im;
    _T_354_re <= _T_353_re;
    _T_354_im <= _T_353_im;
    _T_355_re <= _T_354_re;
    _T_355_im <= _T_354_im;
    _T_356_re <= _T_355_re;
    _T_356_im <= _T_355_im;
    _T_357_re <= _T_356_re;
    _T_357_im <= _T_356_im;
    _T_358_re <= _T_357_re;
    _T_358_im <= _T_357_im;
    _T_359_re <= _T_358_re;
    _T_359_im <= _T_358_im;
    _T_360_re <= _T_359_re;
    _T_360_im <= _T_359_im;
    _T_361_re <= _T_360_re;
    _T_361_im <= _T_360_im;
    _T_362_re <= _T_361_re;
    _T_362_im <= _T_361_im;
    _T_363_re <= _T_362_re;
    _T_363_im <= _T_362_im;
    _T_364_re <= _T_363_re;
    _T_364_im <= _T_363_im;
    _T_365_re <= _T_364_re;
    _T_365_im <= _T_364_im;
    _T_366_re <= _T_365_re;
    _T_366_im <= _T_365_im;
    _T_367_re <= _T_366_re;
    _T_367_im <= _T_366_im;
    _T_368_re <= _T_367_re;
    _T_368_im <= _T_367_im;
    _T_369_re <= _T_368_re;
    _T_369_im <= _T_368_im;
    _T_370_re <= _T_369_re;
    _T_370_im <= _T_369_im;
    _T_371_re <= _T_370_re;
    _T_371_im <= _T_370_im;
    _T_372_re <= _T_371_re;
    _T_372_im <= _T_371_im;
    _T_373_re <= _T_372_re;
    _T_373_im <= _T_372_im;
    _T_374_re <= _T_373_re;
    _T_374_im <= _T_373_im;
    _T_375_re <= _T_374_re;
    _T_375_im <= _T_374_im;
    _T_376_re <= _T_375_re;
    _T_376_im <= _T_375_im;
    _T_377_re <= _T_376_re;
    _T_377_im <= _T_376_im;
    _T_378_re <= _T_377_re;
    _T_378_im <= _T_377_im;
    _T_379_re <= _T_378_re;
    _T_379_im <= _T_378_im;
    _T_380_re <= _T_379_re;
    _T_380_im <= _T_379_im;
    _T_381_re <= _T_380_re;
    _T_381_im <= _T_380_im;
    _T_382_re <= _T_381_re;
    _T_382_im <= _T_381_im;
    _T_383_re <= _T_382_re;
    _T_383_im <= _T_382_im;
    _T_384_re <= _T_383_re;
    _T_384_im <= _T_383_im;
    _T_385_re <= _T_384_re;
    _T_385_im <= _T_384_im;
    _T_386_re <= _T_385_re;
    _T_386_im <= _T_385_im;
    _T_387_re <= _T_386_re;
    _T_387_im <= _T_386_im;
    _T_388_re <= _T_387_re;
    _T_388_im <= _T_387_im;
    _T_389_re <= _T_388_re;
    _T_389_im <= _T_388_im;
    _T_390_re <= _T_389_re;
    _T_390_im <= _T_389_im;
    _T_391_re <= _T_390_re;
    _T_391_im <= _T_390_im;
    _T_392_re <= _T_391_re;
    _T_392_im <= _T_391_im;
    _T_393_re <= _T_392_re;
    _T_393_im <= _T_392_im;
    _T_394_re <= _T_393_re;
    _T_394_im <= _T_393_im;
    _T_395_re <= _T_394_re;
    _T_395_im <= _T_394_im;
    _T_396_re <= _T_395_re;
    _T_396_im <= _T_395_im;
    _T_397_re <= _T_396_re;
    _T_397_im <= _T_396_im;
    _T_398_re <= _T_397_re;
    _T_398_im <= _T_397_im;
    _T_399_re <= _T_398_re;
    _T_399_im <= _T_398_im;
    _T_400_re <= _T_399_re;
    _T_400_im <= _T_399_im;
    _T_401_re <= _T_400_re;
    _T_401_im <= _T_400_im;
    _T_402_re <= _T_401_re;
    _T_402_im <= _T_401_im;
    _T_403_re <= _T_402_re;
    _T_403_im <= _T_402_im;
    _T_404_re <= _T_403_re;
    _T_404_im <= _T_403_im;
    _T_405_re <= _T_404_re;
    _T_405_im <= _T_404_im;
    _T_407_re <= Butterfly_io_out2_re;
    _T_407_im <= Butterfly_io_out2_im;
    _T_408_re <= _T_407_re;
    _T_408_im <= _T_407_im;
    _T_409_re <= _T_408_re;
    _T_409_im <= _T_408_im;
    _T_410_re <= _T_409_re;
    _T_410_im <= _T_409_im;
    _T_411_re <= _T_410_re;
    _T_411_im <= _T_410_im;
    _T_412_re <= _T_411_re;
    _T_412_im <= _T_411_im;
    _T_413_re <= _T_412_re;
    _T_413_im <= _T_412_im;
    _T_414_re <= _T_413_re;
    _T_414_im <= _T_413_im;
    _T_415_re <= _T_414_re;
    _T_415_im <= _T_414_im;
    _T_416_re <= _T_415_re;
    _T_416_im <= _T_415_im;
    _T_417_re <= _T_416_re;
    _T_417_im <= _T_416_im;
    _T_418_re <= _T_417_re;
    _T_418_im <= _T_417_im;
    _T_419_re <= _T_418_re;
    _T_419_im <= _T_418_im;
    _T_420_re <= _T_419_re;
    _T_420_im <= _T_419_im;
    _T_421_re <= _T_420_re;
    _T_421_im <= _T_420_im;
    _T_422_re <= _T_421_re;
    _T_422_im <= _T_421_im;
    _T_423_re <= _T_422_re;
    _T_423_im <= _T_422_im;
    _T_424_re <= _T_423_re;
    _T_424_im <= _T_423_im;
    _T_425_re <= _T_424_re;
    _T_425_im <= _T_424_im;
    _T_426_re <= _T_425_re;
    _T_426_im <= _T_425_im;
    _T_427_re <= _T_426_re;
    _T_427_im <= _T_426_im;
    _T_428_re <= _T_427_re;
    _T_428_im <= _T_427_im;
    _T_429_re <= _T_428_re;
    _T_429_im <= _T_428_im;
    _T_430_re <= _T_429_re;
    _T_430_im <= _T_429_im;
    _T_431_re <= _T_430_re;
    _T_431_im <= _T_430_im;
    _T_432_re <= _T_431_re;
    _T_432_im <= _T_431_im;
    _T_433_re <= _T_432_re;
    _T_433_im <= _T_432_im;
    _T_434_re <= _T_433_re;
    _T_434_im <= _T_433_im;
    _T_435_re <= _T_434_re;
    _T_435_im <= _T_434_im;
    _T_436_re <= _T_435_re;
    _T_436_im <= _T_435_im;
    _T_437_re <= _T_436_re;
    _T_437_im <= _T_436_im;
    _T_438_re <= _T_437_re;
    _T_438_im <= _T_437_im;
    _T_439_re <= _T_438_re;
    _T_439_im <= _T_438_im;
    _T_440_re <= _T_439_re;
    _T_440_im <= _T_439_im;
    _T_441_re <= _T_440_re;
    _T_441_im <= _T_440_im;
    _T_442_re <= _T_441_re;
    _T_442_im <= _T_441_im;
    _T_443_re <= _T_442_re;
    _T_443_im <= _T_442_im;
    _T_444_re <= _T_443_re;
    _T_444_im <= _T_443_im;
    _T_445_re <= _T_444_re;
    _T_445_im <= _T_444_im;
    _T_446_re <= _T_445_re;
    _T_446_im <= _T_445_im;
    _T_447_re <= _T_446_re;
    _T_447_im <= _T_446_im;
    _T_448_re <= _T_447_re;
    _T_448_im <= _T_447_im;
    _T_449_re <= _T_448_re;
    _T_449_im <= _T_448_im;
    _T_450_re <= _T_449_re;
    _T_450_im <= _T_449_im;
    _T_451_re <= _T_450_re;
    _T_451_im <= _T_450_im;
    _T_452_re <= _T_451_re;
    _T_452_im <= _T_451_im;
    _T_453_re <= _T_452_re;
    _T_453_im <= _T_452_im;
    _T_454_re <= _T_453_re;
    _T_454_im <= _T_453_im;
    _T_455_re <= _T_454_re;
    _T_455_im <= _T_454_im;
    _T_456_re <= _T_455_re;
    _T_456_im <= _T_455_im;
    _T_457_re <= _T_456_re;
    _T_457_im <= _T_456_im;
    _T_458_re <= _T_457_re;
    _T_458_im <= _T_457_im;
    _T_459_re <= _T_458_re;
    _T_459_im <= _T_458_im;
    _T_460_re <= _T_459_re;
    _T_460_im <= _T_459_im;
    _T_461_re <= _T_460_re;
    _T_461_im <= _T_460_im;
    _T_462_re <= _T_461_re;
    _T_462_im <= _T_461_im;
    _T_463_re <= _T_462_re;
    _T_463_im <= _T_462_im;
    _T_464_re <= _T_463_re;
    _T_464_im <= _T_463_im;
    _T_465_re <= _T_464_re;
    _T_465_im <= _T_464_im;
    _T_466_re <= _T_465_re;
    _T_466_im <= _T_465_im;
    _T_467_re <= _T_466_re;
    _T_467_im <= _T_466_im;
    _T_468_re <= _T_467_re;
    _T_468_im <= _T_467_im;
    _T_469_re <= _T_468_re;
    _T_469_im <= _T_468_im;
    _T_470_re <= _T_469_re;
    _T_470_im <= _T_469_im;
    _T_471_re <= _T_470_re;
    _T_471_im <= _T_470_im;
    _T_472_re <= _T_471_re;
    _T_472_im <= _T_471_im;
    _T_473_re <= _T_472_re;
    _T_473_im <= _T_472_im;
    _T_474_re <= _T_473_re;
    _T_474_im <= _T_473_im;
    _T_475_re <= _T_474_re;
    _T_475_im <= _T_474_im;
    _T_476_re <= _T_475_re;
    _T_476_im <= _T_475_im;
    _T_477_re <= _T_476_re;
    _T_477_im <= _T_476_im;
    _T_478_re <= _T_477_re;
    _T_478_im <= _T_477_im;
    _T_479_re <= _T_478_re;
    _T_479_im <= _T_478_im;
    _T_480_re <= _T_479_re;
    _T_480_im <= _T_479_im;
    _T_481_re <= _T_480_re;
    _T_481_im <= _T_480_im;
    _T_482_re <= _T_481_re;
    _T_482_im <= _T_481_im;
    _T_483_re <= _T_482_re;
    _T_483_im <= _T_482_im;
    _T_484_re <= _T_483_re;
    _T_484_im <= _T_483_im;
    _T_485_re <= _T_484_re;
    _T_485_im <= _T_484_im;
    _T_486_re <= _T_485_re;
    _T_486_im <= _T_485_im;
    _T_487_re <= _T_486_re;
    _T_487_im <= _T_486_im;
    _T_488_re <= _T_487_re;
    _T_488_im <= _T_487_im;
    _T_489_re <= _T_488_re;
    _T_489_im <= _T_488_im;
    _T_490_re <= _T_489_re;
    _T_490_im <= _T_489_im;
    _T_491_re <= _T_490_re;
    _T_491_im <= _T_490_im;
    _T_492_re <= _T_491_re;
    _T_492_im <= _T_491_im;
    _T_493_re <= _T_492_re;
    _T_493_im <= _T_492_im;
    _T_494_re <= _T_493_re;
    _T_494_im <= _T_493_im;
    _T_495_re <= _T_494_re;
    _T_495_im <= _T_494_im;
    _T_496_re <= _T_495_re;
    _T_496_im <= _T_495_im;
    _T_497_re <= _T_496_re;
    _T_497_im <= _T_496_im;
    _T_498_re <= _T_497_re;
    _T_498_im <= _T_497_im;
    _T_499_re <= _T_498_re;
    _T_499_im <= _T_498_im;
    _T_500_re <= _T_499_re;
    _T_500_im <= _T_499_im;
    _T_501_re <= _T_500_re;
    _T_501_im <= _T_500_im;
    _T_502_re <= _T_501_re;
    _T_502_im <= _T_501_im;
    _T_503_re <= _T_502_re;
    _T_503_im <= _T_502_im;
    _T_504_re <= _T_503_re;
    _T_504_im <= _T_503_im;
    _T_505_re <= _T_504_re;
    _T_505_im <= _T_504_im;
    _T_506_re <= _T_505_re;
    _T_506_im <= _T_505_im;
    _T_507_re <= _T_506_re;
    _T_507_im <= _T_506_im;
    _T_508_re <= _T_507_re;
    _T_508_im <= _T_507_im;
    _T_509_re <= _T_508_re;
    _T_509_im <= _T_508_im;
    _T_510_re <= _T_509_re;
    _T_510_im <= _T_509_im;
    _T_511_re <= _T_510_re;
    _T_511_im <= _T_510_im;
    _T_512_re <= _T_511_re;
    _T_512_im <= _T_511_im;
    _T_513_re <= _T_512_re;
    _T_513_im <= _T_512_im;
    _T_514_re <= _T_513_re;
    _T_514_im <= _T_513_im;
    _T_515_re <= _T_514_re;
    _T_515_im <= _T_514_im;
    _T_516_re <= _T_515_re;
    _T_516_im <= _T_515_im;
    _T_517_re <= _T_516_re;
    _T_517_im <= _T_516_im;
    _T_518_re <= _T_517_re;
    _T_518_im <= _T_517_im;
    _T_519_re <= _T_518_re;
    _T_519_im <= _T_518_im;
    _T_520_re <= _T_519_re;
    _T_520_im <= _T_519_im;
    _T_521_re <= _T_520_re;
    _T_521_im <= _T_520_im;
    _T_522_re <= _T_521_re;
    _T_522_im <= _T_521_im;
    _T_523_re <= _T_522_re;
    _T_523_im <= _T_522_im;
    _T_524_re <= _T_523_re;
    _T_524_im <= _T_523_im;
    _T_525_re <= _T_524_re;
    _T_525_im <= _T_524_im;
    _T_526_re <= _T_525_re;
    _T_526_im <= _T_525_im;
    _T_527_re <= _T_526_re;
    _T_527_im <= _T_526_im;
    _T_528_re <= _T_527_re;
    _T_528_im <= _T_527_im;
    _T_529_re <= _T_528_re;
    _T_529_im <= _T_528_im;
    _T_530_re <= _T_529_re;
    _T_530_im <= _T_529_im;
    _T_531_re <= _T_530_re;
    _T_531_im <= _T_530_im;
    _T_532_re <= _T_531_re;
    _T_532_im <= _T_531_im;
    _T_533_re <= _T_532_re;
    _T_533_im <= _T_532_im;
    _T_534_re <= _T_533_re;
    _T_534_im <= _T_533_im;
    _T_543_re <= Switch_io_out1_re;
    _T_543_im <= Switch_io_out1_im;
    _T_544_re <= _T_543_re;
    _T_544_im <= _T_543_im;
    _T_545_re <= _T_544_re;
    _T_545_im <= _T_544_im;
    _T_546_re <= _T_545_re;
    _T_546_im <= _T_545_im;
    _T_547_re <= _T_546_re;
    _T_547_im <= _T_546_im;
    _T_548_re <= _T_547_re;
    _T_548_im <= _T_547_im;
    _T_549_re <= _T_548_re;
    _T_549_im <= _T_548_im;
    _T_550_re <= _T_549_re;
    _T_550_im <= _T_549_im;
    _T_551_re <= _T_550_re;
    _T_551_im <= _T_550_im;
    _T_552_re <= _T_551_re;
    _T_552_im <= _T_551_im;
    _T_553_re <= _T_552_re;
    _T_553_im <= _T_552_im;
    _T_554_re <= _T_553_re;
    _T_554_im <= _T_553_im;
    _T_555_re <= _T_554_re;
    _T_555_im <= _T_554_im;
    _T_556_re <= _T_555_re;
    _T_556_im <= _T_555_im;
    _T_557_re <= _T_556_re;
    _T_557_im <= _T_556_im;
    _T_558_re <= _T_557_re;
    _T_558_im <= _T_557_im;
    _T_559_re <= _T_558_re;
    _T_559_im <= _T_558_im;
    _T_560_re <= _T_559_re;
    _T_560_im <= _T_559_im;
    _T_561_re <= _T_560_re;
    _T_561_im <= _T_560_im;
    _T_562_re <= _T_561_re;
    _T_562_im <= _T_561_im;
    _T_563_re <= _T_562_re;
    _T_563_im <= _T_562_im;
    _T_564_re <= _T_563_re;
    _T_564_im <= _T_563_im;
    _T_565_re <= _T_564_re;
    _T_565_im <= _T_564_im;
    _T_566_re <= _T_565_re;
    _T_566_im <= _T_565_im;
    _T_567_re <= _T_566_re;
    _T_567_im <= _T_566_im;
    _T_568_re <= _T_567_re;
    _T_568_im <= _T_567_im;
    _T_569_re <= _T_568_re;
    _T_569_im <= _T_568_im;
    _T_570_re <= _T_569_re;
    _T_570_im <= _T_569_im;
    _T_571_re <= _T_570_re;
    _T_571_im <= _T_570_im;
    _T_572_re <= _T_571_re;
    _T_572_im <= _T_571_im;
    _T_573_re <= _T_572_re;
    _T_573_im <= _T_572_im;
    _T_574_re <= _T_573_re;
    _T_574_im <= _T_573_im;
    _T_575_re <= _T_574_re;
    _T_575_im <= _T_574_im;
    _T_576_re <= _T_575_re;
    _T_576_im <= _T_575_im;
    _T_577_re <= _T_576_re;
    _T_577_im <= _T_576_im;
    _T_578_re <= _T_577_re;
    _T_578_im <= _T_577_im;
    _T_579_re <= _T_578_re;
    _T_579_im <= _T_578_im;
    _T_580_re <= _T_579_re;
    _T_580_im <= _T_579_im;
    _T_581_re <= _T_580_re;
    _T_581_im <= _T_580_im;
    _T_582_re <= _T_581_re;
    _T_582_im <= _T_581_im;
    _T_583_re <= _T_582_re;
    _T_583_im <= _T_582_im;
    _T_584_re <= _T_583_re;
    _T_584_im <= _T_583_im;
    _T_585_re <= _T_584_re;
    _T_585_im <= _T_584_im;
    _T_586_re <= _T_585_re;
    _T_586_im <= _T_585_im;
    _T_587_re <= _T_586_re;
    _T_587_im <= _T_586_im;
    _T_588_re <= _T_587_re;
    _T_588_im <= _T_587_im;
    _T_589_re <= _T_588_re;
    _T_589_im <= _T_588_im;
    _T_590_re <= _T_589_re;
    _T_590_im <= _T_589_im;
    _T_591_re <= _T_590_re;
    _T_591_im <= _T_590_im;
    _T_592_re <= _T_591_re;
    _T_592_im <= _T_591_im;
    _T_593_re <= _T_592_re;
    _T_593_im <= _T_592_im;
    _T_594_re <= _T_593_re;
    _T_594_im <= _T_593_im;
    _T_595_re <= _T_594_re;
    _T_595_im <= _T_594_im;
    _T_596_re <= _T_595_re;
    _T_596_im <= _T_595_im;
    _T_597_re <= _T_596_re;
    _T_597_im <= _T_596_im;
    _T_598_re <= _T_597_re;
    _T_598_im <= _T_597_im;
    _T_599_re <= _T_598_re;
    _T_599_im <= _T_598_im;
    _T_600_re <= _T_599_re;
    _T_600_im <= _T_599_im;
    _T_601_re <= _T_600_re;
    _T_601_im <= _T_600_im;
    _T_602_re <= _T_601_re;
    _T_602_im <= _T_601_im;
    _T_603_re <= _T_602_re;
    _T_603_im <= _T_602_im;
    _T_604_re <= _T_603_re;
    _T_604_im <= _T_603_im;
    _T_605_re <= _T_604_re;
    _T_605_im <= _T_604_im;
    _T_606_re <= _T_605_re;
    _T_606_im <= _T_605_im;
    _T_607_re <= _T_606_re;
    _T_607_im <= _T_606_im;
    _T_608_re <= _T_607_re;
    _T_608_im <= _T_607_im;
    _T_609_re <= _T_608_re;
    _T_609_im <= _T_608_im;
    _T_610_re <= _T_609_re;
    _T_610_im <= _T_609_im;
    _T_611_re <= _T_610_re;
    _T_611_im <= _T_610_im;
    _T_612_re <= _T_611_re;
    _T_612_im <= _T_611_im;
    _T_613_re <= _T_612_re;
    _T_613_im <= _T_612_im;
    _T_614_re <= _T_613_re;
    _T_614_im <= _T_613_im;
    _T_615_re <= _T_614_re;
    _T_615_im <= _T_614_im;
    _T_616_re <= _T_615_re;
    _T_616_im <= _T_615_im;
    _T_617_re <= _T_616_re;
    _T_617_im <= _T_616_im;
    _T_618_re <= _T_617_re;
    _T_618_im <= _T_617_im;
    _T_619_re <= _T_618_re;
    _T_619_im <= _T_618_im;
    _T_620_re <= _T_619_re;
    _T_620_im <= _T_619_im;
    _T_621_re <= _T_620_re;
    _T_621_im <= _T_620_im;
    _T_622_re <= _T_621_re;
    _T_622_im <= _T_621_im;
    _T_623_re <= _T_622_re;
    _T_623_im <= _T_622_im;
    _T_624_re <= _T_623_re;
    _T_624_im <= _T_623_im;
    _T_625_re <= _T_624_re;
    _T_625_im <= _T_624_im;
    _T_626_re <= _T_625_re;
    _T_626_im <= _T_625_im;
    _T_627_re <= _T_626_re;
    _T_627_im <= _T_626_im;
    _T_628_re <= _T_627_re;
    _T_628_im <= _T_627_im;
    _T_629_re <= _T_628_re;
    _T_629_im <= _T_628_im;
    _T_630_re <= _T_629_re;
    _T_630_im <= _T_629_im;
    _T_631_re <= _T_630_re;
    _T_631_im <= _T_630_im;
    _T_632_re <= _T_631_re;
    _T_632_im <= _T_631_im;
    _T_633_re <= _T_632_re;
    _T_633_im <= _T_632_im;
    _T_634_re <= _T_633_re;
    _T_634_im <= _T_633_im;
    _T_635_re <= _T_634_re;
    _T_635_im <= _T_634_im;
    _T_636_re <= _T_635_re;
    _T_636_im <= _T_635_im;
    _T_637_re <= _T_636_re;
    _T_637_im <= _T_636_im;
    _T_638_re <= _T_637_re;
    _T_638_im <= _T_637_im;
    _T_639_re <= _T_638_re;
    _T_639_im <= _T_638_im;
    _T_640_re <= _T_639_re;
    _T_640_im <= _T_639_im;
    _T_641_re <= _T_640_re;
    _T_641_im <= _T_640_im;
    _T_642_re <= _T_641_re;
    _T_642_im <= _T_641_im;
    _T_643_re <= _T_642_re;
    _T_643_im <= _T_642_im;
    _T_644_re <= _T_643_re;
    _T_644_im <= _T_643_im;
    _T_645_re <= _T_644_re;
    _T_645_im <= _T_644_im;
    _T_646_re <= _T_645_re;
    _T_646_im <= _T_645_im;
    _T_647_re <= _T_646_re;
    _T_647_im <= _T_646_im;
    _T_648_re <= _T_647_re;
    _T_648_im <= _T_647_im;
    _T_649_re <= _T_648_re;
    _T_649_im <= _T_648_im;
    _T_650_re <= _T_649_re;
    _T_650_im <= _T_649_im;
    _T_651_re <= _T_650_re;
    _T_651_im <= _T_650_im;
    _T_652_re <= _T_651_re;
    _T_652_im <= _T_651_im;
    _T_653_re <= _T_652_re;
    _T_653_im <= _T_652_im;
    _T_654_re <= _T_653_re;
    _T_654_im <= _T_653_im;
    _T_655_re <= _T_654_re;
    _T_655_im <= _T_654_im;
    _T_656_re <= _T_655_re;
    _T_656_im <= _T_655_im;
    _T_657_re <= _T_656_re;
    _T_657_im <= _T_656_im;
    _T_658_re <= _T_657_re;
    _T_658_im <= _T_657_im;
    _T_659_re <= _T_658_re;
    _T_659_im <= _T_658_im;
    _T_660_re <= _T_659_re;
    _T_660_im <= _T_659_im;
    _T_661_re <= _T_660_re;
    _T_661_im <= _T_660_im;
    _T_662_re <= _T_661_re;
    _T_662_im <= _T_661_im;
    _T_663_re <= _T_662_re;
    _T_663_im <= _T_662_im;
    _T_664_re <= _T_663_re;
    _T_664_im <= _T_663_im;
    _T_665_re <= _T_664_re;
    _T_665_im <= _T_664_im;
    _T_666_re <= _T_665_re;
    _T_666_im <= _T_665_im;
    _T_667_re <= _T_666_re;
    _T_667_im <= _T_666_im;
    _T_668_re <= _T_667_re;
    _T_668_im <= _T_667_im;
    _T_669_re <= _T_668_re;
    _T_669_im <= _T_668_im;
    _T_670_re <= _T_669_re;
    _T_670_im <= _T_669_im;
    _T_672_re <= Butterfly_1_io_out2_re;
    _T_672_im <= Butterfly_1_io_out2_im;
    _T_673_re <= _T_672_re;
    _T_673_im <= _T_672_im;
    _T_674_re <= _T_673_re;
    _T_674_im <= _T_673_im;
    _T_675_re <= _T_674_re;
    _T_675_im <= _T_674_im;
    _T_676_re <= _T_675_re;
    _T_676_im <= _T_675_im;
    _T_677_re <= _T_676_re;
    _T_677_im <= _T_676_im;
    _T_678_re <= _T_677_re;
    _T_678_im <= _T_677_im;
    _T_679_re <= _T_678_re;
    _T_679_im <= _T_678_im;
    _T_680_re <= _T_679_re;
    _T_680_im <= _T_679_im;
    _T_681_re <= _T_680_re;
    _T_681_im <= _T_680_im;
    _T_682_re <= _T_681_re;
    _T_682_im <= _T_681_im;
    _T_683_re <= _T_682_re;
    _T_683_im <= _T_682_im;
    _T_684_re <= _T_683_re;
    _T_684_im <= _T_683_im;
    _T_685_re <= _T_684_re;
    _T_685_im <= _T_684_im;
    _T_686_re <= _T_685_re;
    _T_686_im <= _T_685_im;
    _T_687_re <= _T_686_re;
    _T_687_im <= _T_686_im;
    _T_688_re <= _T_687_re;
    _T_688_im <= _T_687_im;
    _T_689_re <= _T_688_re;
    _T_689_im <= _T_688_im;
    _T_690_re <= _T_689_re;
    _T_690_im <= _T_689_im;
    _T_691_re <= _T_690_re;
    _T_691_im <= _T_690_im;
    _T_692_re <= _T_691_re;
    _T_692_im <= _T_691_im;
    _T_693_re <= _T_692_re;
    _T_693_im <= _T_692_im;
    _T_694_re <= _T_693_re;
    _T_694_im <= _T_693_im;
    _T_695_re <= _T_694_re;
    _T_695_im <= _T_694_im;
    _T_696_re <= _T_695_re;
    _T_696_im <= _T_695_im;
    _T_697_re <= _T_696_re;
    _T_697_im <= _T_696_im;
    _T_698_re <= _T_697_re;
    _T_698_im <= _T_697_im;
    _T_699_re <= _T_698_re;
    _T_699_im <= _T_698_im;
    _T_700_re <= _T_699_re;
    _T_700_im <= _T_699_im;
    _T_701_re <= _T_700_re;
    _T_701_im <= _T_700_im;
    _T_702_re <= _T_701_re;
    _T_702_im <= _T_701_im;
    _T_703_re <= _T_702_re;
    _T_703_im <= _T_702_im;
    _T_704_re <= _T_703_re;
    _T_704_im <= _T_703_im;
    _T_705_re <= _T_704_re;
    _T_705_im <= _T_704_im;
    _T_706_re <= _T_705_re;
    _T_706_im <= _T_705_im;
    _T_707_re <= _T_706_re;
    _T_707_im <= _T_706_im;
    _T_708_re <= _T_707_re;
    _T_708_im <= _T_707_im;
    _T_709_re <= _T_708_re;
    _T_709_im <= _T_708_im;
    _T_710_re <= _T_709_re;
    _T_710_im <= _T_709_im;
    _T_711_re <= _T_710_re;
    _T_711_im <= _T_710_im;
    _T_712_re <= _T_711_re;
    _T_712_im <= _T_711_im;
    _T_713_re <= _T_712_re;
    _T_713_im <= _T_712_im;
    _T_714_re <= _T_713_re;
    _T_714_im <= _T_713_im;
    _T_715_re <= _T_714_re;
    _T_715_im <= _T_714_im;
    _T_716_re <= _T_715_re;
    _T_716_im <= _T_715_im;
    _T_717_re <= _T_716_re;
    _T_717_im <= _T_716_im;
    _T_718_re <= _T_717_re;
    _T_718_im <= _T_717_im;
    _T_719_re <= _T_718_re;
    _T_719_im <= _T_718_im;
    _T_720_re <= _T_719_re;
    _T_720_im <= _T_719_im;
    _T_721_re <= _T_720_re;
    _T_721_im <= _T_720_im;
    _T_722_re <= _T_721_re;
    _T_722_im <= _T_721_im;
    _T_723_re <= _T_722_re;
    _T_723_im <= _T_722_im;
    _T_724_re <= _T_723_re;
    _T_724_im <= _T_723_im;
    _T_725_re <= _T_724_re;
    _T_725_im <= _T_724_im;
    _T_726_re <= _T_725_re;
    _T_726_im <= _T_725_im;
    _T_727_re <= _T_726_re;
    _T_727_im <= _T_726_im;
    _T_728_re <= _T_727_re;
    _T_728_im <= _T_727_im;
    _T_729_re <= _T_728_re;
    _T_729_im <= _T_728_im;
    _T_730_re <= _T_729_re;
    _T_730_im <= _T_729_im;
    _T_731_re <= _T_730_re;
    _T_731_im <= _T_730_im;
    _T_732_re <= _T_731_re;
    _T_732_im <= _T_731_im;
    _T_733_re <= _T_732_re;
    _T_733_im <= _T_732_im;
    _T_734_re <= _T_733_re;
    _T_734_im <= _T_733_im;
    _T_735_re <= _T_734_re;
    _T_735_im <= _T_734_im;
    _T_744_re <= Switch_1_io_out1_re;
    _T_744_im <= Switch_1_io_out1_im;
    _T_745_re <= _T_744_re;
    _T_745_im <= _T_744_im;
    _T_746_re <= _T_745_re;
    _T_746_im <= _T_745_im;
    _T_747_re <= _T_746_re;
    _T_747_im <= _T_746_im;
    _T_748_re <= _T_747_re;
    _T_748_im <= _T_747_im;
    _T_749_re <= _T_748_re;
    _T_749_im <= _T_748_im;
    _T_750_re <= _T_749_re;
    _T_750_im <= _T_749_im;
    _T_751_re <= _T_750_re;
    _T_751_im <= _T_750_im;
    _T_752_re <= _T_751_re;
    _T_752_im <= _T_751_im;
    _T_753_re <= _T_752_re;
    _T_753_im <= _T_752_im;
    _T_754_re <= _T_753_re;
    _T_754_im <= _T_753_im;
    _T_755_re <= _T_754_re;
    _T_755_im <= _T_754_im;
    _T_756_re <= _T_755_re;
    _T_756_im <= _T_755_im;
    _T_757_re <= _T_756_re;
    _T_757_im <= _T_756_im;
    _T_758_re <= _T_757_re;
    _T_758_im <= _T_757_im;
    _T_759_re <= _T_758_re;
    _T_759_im <= _T_758_im;
    _T_760_re <= _T_759_re;
    _T_760_im <= _T_759_im;
    _T_761_re <= _T_760_re;
    _T_761_im <= _T_760_im;
    _T_762_re <= _T_761_re;
    _T_762_im <= _T_761_im;
    _T_763_re <= _T_762_re;
    _T_763_im <= _T_762_im;
    _T_764_re <= _T_763_re;
    _T_764_im <= _T_763_im;
    _T_765_re <= _T_764_re;
    _T_765_im <= _T_764_im;
    _T_766_re <= _T_765_re;
    _T_766_im <= _T_765_im;
    _T_767_re <= _T_766_re;
    _T_767_im <= _T_766_im;
    _T_768_re <= _T_767_re;
    _T_768_im <= _T_767_im;
    _T_769_re <= _T_768_re;
    _T_769_im <= _T_768_im;
    _T_770_re <= _T_769_re;
    _T_770_im <= _T_769_im;
    _T_771_re <= _T_770_re;
    _T_771_im <= _T_770_im;
    _T_772_re <= _T_771_re;
    _T_772_im <= _T_771_im;
    _T_773_re <= _T_772_re;
    _T_773_im <= _T_772_im;
    _T_774_re <= _T_773_re;
    _T_774_im <= _T_773_im;
    _T_775_re <= _T_774_re;
    _T_775_im <= _T_774_im;
    _T_776_re <= _T_775_re;
    _T_776_im <= _T_775_im;
    _T_777_re <= _T_776_re;
    _T_777_im <= _T_776_im;
    _T_778_re <= _T_777_re;
    _T_778_im <= _T_777_im;
    _T_779_re <= _T_778_re;
    _T_779_im <= _T_778_im;
    _T_780_re <= _T_779_re;
    _T_780_im <= _T_779_im;
    _T_781_re <= _T_780_re;
    _T_781_im <= _T_780_im;
    _T_782_re <= _T_781_re;
    _T_782_im <= _T_781_im;
    _T_783_re <= _T_782_re;
    _T_783_im <= _T_782_im;
    _T_784_re <= _T_783_re;
    _T_784_im <= _T_783_im;
    _T_785_re <= _T_784_re;
    _T_785_im <= _T_784_im;
    _T_786_re <= _T_785_re;
    _T_786_im <= _T_785_im;
    _T_787_re <= _T_786_re;
    _T_787_im <= _T_786_im;
    _T_788_re <= _T_787_re;
    _T_788_im <= _T_787_im;
    _T_789_re <= _T_788_re;
    _T_789_im <= _T_788_im;
    _T_790_re <= _T_789_re;
    _T_790_im <= _T_789_im;
    _T_791_re <= _T_790_re;
    _T_791_im <= _T_790_im;
    _T_792_re <= _T_791_re;
    _T_792_im <= _T_791_im;
    _T_793_re <= _T_792_re;
    _T_793_im <= _T_792_im;
    _T_794_re <= _T_793_re;
    _T_794_im <= _T_793_im;
    _T_795_re <= _T_794_re;
    _T_795_im <= _T_794_im;
    _T_796_re <= _T_795_re;
    _T_796_im <= _T_795_im;
    _T_797_re <= _T_796_re;
    _T_797_im <= _T_796_im;
    _T_798_re <= _T_797_re;
    _T_798_im <= _T_797_im;
    _T_799_re <= _T_798_re;
    _T_799_im <= _T_798_im;
    _T_800_re <= _T_799_re;
    _T_800_im <= _T_799_im;
    _T_801_re <= _T_800_re;
    _T_801_im <= _T_800_im;
    _T_802_re <= _T_801_re;
    _T_802_im <= _T_801_im;
    _T_803_re <= _T_802_re;
    _T_803_im <= _T_802_im;
    _T_804_re <= _T_803_re;
    _T_804_im <= _T_803_im;
    _T_805_re <= _T_804_re;
    _T_805_im <= _T_804_im;
    _T_806_re <= _T_805_re;
    _T_806_im <= _T_805_im;
    _T_807_re <= _T_806_re;
    _T_807_im <= _T_806_im;
    _T_809_re <= Butterfly_2_io_out2_re;
    _T_809_im <= Butterfly_2_io_out2_im;
    _T_810_re <= _T_809_re;
    _T_810_im <= _T_809_im;
    _T_811_re <= _T_810_re;
    _T_811_im <= _T_810_im;
    _T_812_re <= _T_811_re;
    _T_812_im <= _T_811_im;
    _T_813_re <= _T_812_re;
    _T_813_im <= _T_812_im;
    _T_814_re <= _T_813_re;
    _T_814_im <= _T_813_im;
    _T_815_re <= _T_814_re;
    _T_815_im <= _T_814_im;
    _T_816_re <= _T_815_re;
    _T_816_im <= _T_815_im;
    _T_817_re <= _T_816_re;
    _T_817_im <= _T_816_im;
    _T_818_re <= _T_817_re;
    _T_818_im <= _T_817_im;
    _T_819_re <= _T_818_re;
    _T_819_im <= _T_818_im;
    _T_820_re <= _T_819_re;
    _T_820_im <= _T_819_im;
    _T_821_re <= _T_820_re;
    _T_821_im <= _T_820_im;
    _T_822_re <= _T_821_re;
    _T_822_im <= _T_821_im;
    _T_823_re <= _T_822_re;
    _T_823_im <= _T_822_im;
    _T_824_re <= _T_823_re;
    _T_824_im <= _T_823_im;
    _T_825_re <= _T_824_re;
    _T_825_im <= _T_824_im;
    _T_826_re <= _T_825_re;
    _T_826_im <= _T_825_im;
    _T_827_re <= _T_826_re;
    _T_827_im <= _T_826_im;
    _T_828_re <= _T_827_re;
    _T_828_im <= _T_827_im;
    _T_829_re <= _T_828_re;
    _T_829_im <= _T_828_im;
    _T_830_re <= _T_829_re;
    _T_830_im <= _T_829_im;
    _T_831_re <= _T_830_re;
    _T_831_im <= _T_830_im;
    _T_832_re <= _T_831_re;
    _T_832_im <= _T_831_im;
    _T_833_re <= _T_832_re;
    _T_833_im <= _T_832_im;
    _T_834_re <= _T_833_re;
    _T_834_im <= _T_833_im;
    _T_835_re <= _T_834_re;
    _T_835_im <= _T_834_im;
    _T_836_re <= _T_835_re;
    _T_836_im <= _T_835_im;
    _T_837_re <= _T_836_re;
    _T_837_im <= _T_836_im;
    _T_838_re <= _T_837_re;
    _T_838_im <= _T_837_im;
    _T_839_re <= _T_838_re;
    _T_839_im <= _T_838_im;
    _T_840_re <= _T_839_re;
    _T_840_im <= _T_839_im;
    _T_849_re <= Switch_2_io_out1_re;
    _T_849_im <= Switch_2_io_out1_im;
    _T_850_re <= _T_849_re;
    _T_850_im <= _T_849_im;
    _T_851_re <= _T_850_re;
    _T_851_im <= _T_850_im;
    _T_852_re <= _T_851_re;
    _T_852_im <= _T_851_im;
    _T_853_re <= _T_852_re;
    _T_853_im <= _T_852_im;
    _T_854_re <= _T_853_re;
    _T_854_im <= _T_853_im;
    _T_855_re <= _T_854_re;
    _T_855_im <= _T_854_im;
    _T_856_re <= _T_855_re;
    _T_856_im <= _T_855_im;
    _T_857_re <= _T_856_re;
    _T_857_im <= _T_856_im;
    _T_858_re <= _T_857_re;
    _T_858_im <= _T_857_im;
    _T_859_re <= _T_858_re;
    _T_859_im <= _T_858_im;
    _T_860_re <= _T_859_re;
    _T_860_im <= _T_859_im;
    _T_861_re <= _T_860_re;
    _T_861_im <= _T_860_im;
    _T_862_re <= _T_861_re;
    _T_862_im <= _T_861_im;
    _T_863_re <= _T_862_re;
    _T_863_im <= _T_862_im;
    _T_864_re <= _T_863_re;
    _T_864_im <= _T_863_im;
    _T_865_re <= _T_864_re;
    _T_865_im <= _T_864_im;
    _T_866_re <= _T_865_re;
    _T_866_im <= _T_865_im;
    _T_867_re <= _T_866_re;
    _T_867_im <= _T_866_im;
    _T_868_re <= _T_867_re;
    _T_868_im <= _T_867_im;
    _T_869_re <= _T_868_re;
    _T_869_im <= _T_868_im;
    _T_870_re <= _T_869_re;
    _T_870_im <= _T_869_im;
    _T_871_re <= _T_870_re;
    _T_871_im <= _T_870_im;
    _T_872_re <= _T_871_re;
    _T_872_im <= _T_871_im;
    _T_873_re <= _T_872_re;
    _T_873_im <= _T_872_im;
    _T_874_re <= _T_873_re;
    _T_874_im <= _T_873_im;
    _T_875_re <= _T_874_re;
    _T_875_im <= _T_874_im;
    _T_876_re <= _T_875_re;
    _T_876_im <= _T_875_im;
    _T_877_re <= _T_876_re;
    _T_877_im <= _T_876_im;
    _T_878_re <= _T_877_re;
    _T_878_im <= _T_877_im;
    _T_879_re <= _T_878_re;
    _T_879_im <= _T_878_im;
    _T_880_re <= _T_879_re;
    _T_880_im <= _T_879_im;
    _T_882_re <= Butterfly_3_io_out2_re;
    _T_882_im <= Butterfly_3_io_out2_im;
    _T_883_re <= _T_882_re;
    _T_883_im <= _T_882_im;
    _T_884_re <= _T_883_re;
    _T_884_im <= _T_883_im;
    _T_885_re <= _T_884_re;
    _T_885_im <= _T_884_im;
    _T_886_re <= _T_885_re;
    _T_886_im <= _T_885_im;
    _T_887_re <= _T_886_re;
    _T_887_im <= _T_886_im;
    _T_888_re <= _T_887_re;
    _T_888_im <= _T_887_im;
    _T_889_re <= _T_888_re;
    _T_889_im <= _T_888_im;
    _T_890_re <= _T_889_re;
    _T_890_im <= _T_889_im;
    _T_891_re <= _T_890_re;
    _T_891_im <= _T_890_im;
    _T_892_re <= _T_891_re;
    _T_892_im <= _T_891_im;
    _T_893_re <= _T_892_re;
    _T_893_im <= _T_892_im;
    _T_894_re <= _T_893_re;
    _T_894_im <= _T_893_im;
    _T_895_re <= _T_894_re;
    _T_895_im <= _T_894_im;
    _T_896_re <= _T_895_re;
    _T_896_im <= _T_895_im;
    _T_897_re <= _T_896_re;
    _T_897_im <= _T_896_im;
    _T_906_re <= Switch_3_io_out1_re;
    _T_906_im <= Switch_3_io_out1_im;
    _T_907_re <= _T_906_re;
    _T_907_im <= _T_906_im;
    _T_908_re <= _T_907_re;
    _T_908_im <= _T_907_im;
    _T_909_re <= _T_908_re;
    _T_909_im <= _T_908_im;
    _T_910_re <= _T_909_re;
    _T_910_im <= _T_909_im;
    _T_911_re <= _T_910_re;
    _T_911_im <= _T_910_im;
    _T_912_re <= _T_911_re;
    _T_912_im <= _T_911_im;
    _T_913_re <= _T_912_re;
    _T_913_im <= _T_912_im;
    _T_914_re <= _T_913_re;
    _T_914_im <= _T_913_im;
    _T_915_re <= _T_914_re;
    _T_915_im <= _T_914_im;
    _T_916_re <= _T_915_re;
    _T_916_im <= _T_915_im;
    _T_917_re <= _T_916_re;
    _T_917_im <= _T_916_im;
    _T_918_re <= _T_917_re;
    _T_918_im <= _T_917_im;
    _T_919_re <= _T_918_re;
    _T_919_im <= _T_918_im;
    _T_920_re <= _T_919_re;
    _T_920_im <= _T_919_im;
    _T_921_re <= _T_920_re;
    _T_921_im <= _T_920_im;
    _T_923_re <= Butterfly_4_io_out2_re;
    _T_923_im <= Butterfly_4_io_out2_im;
    _T_924_re <= _T_923_re;
    _T_924_im <= _T_923_im;
    _T_925_re <= _T_924_re;
    _T_925_im <= _T_924_im;
    _T_926_re <= _T_925_re;
    _T_926_im <= _T_925_im;
    _T_927_re <= _T_926_re;
    _T_927_im <= _T_926_im;
    _T_928_re <= _T_927_re;
    _T_928_im <= _T_927_im;
    _T_929_re <= _T_928_re;
    _T_929_im <= _T_928_im;
    _T_930_re <= _T_929_re;
    _T_930_im <= _T_929_im;
    _T_939_re <= Switch_4_io_out1_re;
    _T_939_im <= Switch_4_io_out1_im;
    _T_940_re <= _T_939_re;
    _T_940_im <= _T_939_im;
    _T_941_re <= _T_940_re;
    _T_941_im <= _T_940_im;
    _T_942_re <= _T_941_re;
    _T_942_im <= _T_941_im;
    _T_943_re <= _T_942_re;
    _T_943_im <= _T_942_im;
    _T_944_re <= _T_943_re;
    _T_944_im <= _T_943_im;
    _T_945_re <= _T_944_re;
    _T_945_im <= _T_944_im;
    _T_946_re <= _T_945_re;
    _T_946_im <= _T_945_im;
    _T_948_re <= Butterfly_5_io_out2_re;
    _T_948_im <= Butterfly_5_io_out2_im;
    _T_949_re <= _T_948_re;
    _T_949_im <= _T_948_im;
    _T_950_re <= _T_949_re;
    _T_950_im <= _T_949_im;
    _T_951_re <= _T_950_re;
    _T_951_im <= _T_950_im;
    _T_960_re <= Switch_5_io_out1_re;
    _T_960_im <= Switch_5_io_out1_im;
    _T_961_re <= _T_960_re;
    _T_961_im <= _T_960_im;
    _T_962_re <= _T_961_re;
    _T_962_im <= _T_961_im;
    _T_963_re <= _T_962_re;
    _T_963_im <= _T_962_im;
    _T_965_re <= Butterfly_6_io_out2_re;
    _T_965_im <= Butterfly_6_io_out2_im;
    _T_966_re <= _T_965_re;
    _T_966_im <= _T_965_im;
    _T_975_re <= Switch_6_io_out1_re;
    _T_975_im <= Switch_6_io_out1_im;
    _T_976_re <= _T_975_re;
    _T_976_im <= _T_975_im;
    _T_978_re <= Butterfly_7_io_out2_re;
    _T_978_im <= Butterfly_7_io_out2_im;
    out1D1_re <= Switch_7_io_out1_re;
    out1D1_im <= Switch_7_io_out1_im;
    _T_985_re <= ComplexAdd_io_res_re;
    _T_985_im <= ComplexAdd_io_res_im;
    _T_986_re <= ComplexSub_io_res_re;
    _T_986_im <= ComplexSub_io_res_im;
    _T_987 <= io_din_valid;
    _T_988 <= _T_987;
    _T_989 <= _T_988;
    _T_990 <= _T_989;
    _T_991 <= _T_990;
    _T_992 <= _T_991;
    _T_993 <= _T_992;
    _T_994 <= _T_993;
    _T_995 <= _T_994;
    _T_996 <= _T_995;
    _T_997 <= _T_996;
    _T_998 <= _T_997;
    _T_999 <= _T_998;
    _T_1000 <= _T_999;
    _T_1001 <= _T_1000;
    _T_1002 <= _T_1001;
    _T_1003 <= _T_1002;
    _T_1004 <= _T_1003;
    _T_1005 <= _T_1004;
    _T_1006 <= _T_1005;
    _T_1007 <= _T_1006;
    _T_1008 <= _T_1007;
    _T_1009 <= _T_1008;
    _T_1010 <= _T_1009;
    _T_1011 <= _T_1010;
    _T_1012 <= _T_1011;
    _T_1013 <= _T_1012;
    _T_1014 <= _T_1013;
    _T_1015 <= _T_1014;
    _T_1016 <= _T_1015;
    _T_1017 <= _T_1016;
    _T_1018 <= _T_1017;
    _T_1019 <= _T_1018;
    _T_1020 <= _T_1019;
    _T_1021 <= _T_1020;
    _T_1022 <= _T_1021;
    _T_1023 <= _T_1022;
    _T_1024 <= _T_1023;
    _T_1025 <= _T_1024;
    _T_1026 <= _T_1025;
    _T_1027 <= _T_1026;
    _T_1028 <= _T_1027;
    _T_1029 <= _T_1028;
    _T_1030 <= _T_1029;
    _T_1031 <= _T_1030;
    _T_1032 <= _T_1031;
    _T_1033 <= _T_1032;
    _T_1034 <= _T_1033;
    _T_1035 <= _T_1034;
    _T_1036 <= _T_1035;
    _T_1037 <= _T_1036;
    _T_1038 <= _T_1037;
    _T_1039 <= _T_1038;
    _T_1040 <= _T_1039;
    _T_1041 <= _T_1040;
    _T_1042 <= _T_1041;
    _T_1043 <= _T_1042;
    _T_1044 <= _T_1043;
    _T_1045 <= _T_1044;
    _T_1046 <= _T_1045;
    _T_1047 <= _T_1046;
    _T_1048 <= _T_1047;
    _T_1049 <= _T_1048;
    _T_1050 <= _T_1049;
    _T_1051 <= _T_1050;
    _T_1052 <= _T_1051;
    _T_1053 <= _T_1052;
    _T_1054 <= _T_1053;
    _T_1055 <= _T_1054;
    _T_1056 <= _T_1055;
    _T_1057 <= _T_1056;
    _T_1058 <= _T_1057;
    _T_1059 <= _T_1058;
    _T_1060 <= _T_1059;
    _T_1061 <= _T_1060;
    _T_1062 <= _T_1061;
    _T_1063 <= _T_1062;
    _T_1064 <= _T_1063;
    _T_1065 <= _T_1064;
    _T_1066 <= _T_1065;
    _T_1067 <= _T_1066;
    _T_1068 <= _T_1067;
    _T_1069 <= _T_1068;
    _T_1070 <= _T_1069;
    _T_1071 <= _T_1070;
    _T_1072 <= _T_1071;
    _T_1073 <= _T_1072;
    _T_1074 <= _T_1073;
    _T_1075 <= _T_1074;
    _T_1076 <= _T_1075;
    _T_1077 <= _T_1076;
    _T_1078 <= _T_1077;
    _T_1079 <= _T_1078;
    _T_1080 <= _T_1079;
    _T_1081 <= _T_1080;
    _T_1082 <= _T_1081;
    _T_1083 <= _T_1082;
    _T_1084 <= _T_1083;
    _T_1085 <= _T_1084;
    _T_1086 <= _T_1085;
    _T_1087 <= _T_1086;
    _T_1088 <= _T_1087;
    _T_1089 <= _T_1088;
    _T_1090 <= _T_1089;
    _T_1091 <= _T_1090;
    _T_1092 <= _T_1091;
    _T_1093 <= _T_1092;
    _T_1094 <= _T_1093;
    _T_1095 <= _T_1094;
    _T_1096 <= _T_1095;
    _T_1097 <= _T_1096;
    _T_1098 <= _T_1097;
    _T_1099 <= _T_1098;
    _T_1100 <= _T_1099;
    _T_1101 <= _T_1100;
    _T_1102 <= _T_1101;
    _T_1103 <= _T_1102;
    _T_1104 <= _T_1103;
    _T_1105 <= _T_1104;
    _T_1106 <= _T_1105;
    _T_1107 <= _T_1106;
    _T_1108 <= _T_1107;
    _T_1109 <= _T_1108;
    _T_1110 <= _T_1109;
    _T_1111 <= _T_1110;
    _T_1112 <= _T_1111;
    _T_1113 <= _T_1112;
    _T_1114 <= _T_1113;
    _T_1115 <= _T_1114;
    _T_1116 <= _T_1115;
    _T_1117 <= _T_1116;
    _T_1118 <= _T_1117;
    _T_1119 <= _T_1118;
    _T_1120 <= _T_1119;
    _T_1121 <= _T_1120;
    _T_1122 <= _T_1121;
    _T_1123 <= _T_1122;
    _T_1124 <= _T_1123;
    _T_1125 <= _T_1124;
    _T_1126 <= _T_1125;
    _T_1127 <= _T_1126;
    _T_1128 <= _T_1127;
    _T_1129 <= _T_1128;
    _T_1130 <= _T_1129;
    _T_1131 <= _T_1130;
    _T_1132 <= _T_1131;
    _T_1133 <= _T_1132;
    _T_1134 <= _T_1133;
    _T_1135 <= _T_1134;
    _T_1136 <= _T_1135;
    _T_1137 <= _T_1136;
    _T_1138 <= _T_1137;
    _T_1139 <= _T_1138;
    _T_1140 <= _T_1139;
    _T_1141 <= _T_1140;
    _T_1142 <= _T_1141;
    _T_1143 <= _T_1142;
    _T_1144 <= _T_1143;
    _T_1145 <= _T_1144;
    _T_1146 <= _T_1145;
    _T_1147 <= _T_1146;
    _T_1148 <= _T_1147;
    _T_1149 <= _T_1148;
    _T_1150 <= _T_1149;
    _T_1151 <= _T_1150;
    _T_1152 <= _T_1151;
    _T_1153 <= _T_1152;
    _T_1154 <= _T_1153;
    _T_1155 <= _T_1154;
    _T_1156 <= _T_1155;
    _T_1157 <= _T_1156;
    _T_1158 <= _T_1157;
    _T_1159 <= _T_1158;
    _T_1160 <= _T_1159;
    _T_1161 <= _T_1160;
    _T_1162 <= _T_1161;
    _T_1163 <= _T_1162;
    _T_1164 <= _T_1163;
    _T_1165 <= _T_1164;
    _T_1166 <= _T_1165;
    _T_1167 <= _T_1166;
    _T_1168 <= _T_1167;
    _T_1169 <= _T_1168;
    _T_1170 <= _T_1169;
    _T_1171 <= _T_1170;
    _T_1172 <= _T_1171;
    _T_1173 <= _T_1172;
    _T_1174 <= _T_1173;
    _T_1175 <= _T_1174;
    _T_1176 <= _T_1175;
    _T_1177 <= _T_1176;
    _T_1178 <= _T_1177;
    _T_1179 <= _T_1178;
    _T_1180 <= _T_1179;
    _T_1181 <= _T_1180;
    _T_1182 <= _T_1181;
    _T_1183 <= _T_1182;
    _T_1184 <= _T_1183;
    _T_1185 <= _T_1184;
    _T_1186 <= _T_1185;
    _T_1187 <= _T_1186;
    _T_1188 <= _T_1187;
    _T_1189 <= _T_1188;
    _T_1190 <= _T_1189;
    _T_1191 <= _T_1190;
    _T_1192 <= _T_1191;
    _T_1193 <= _T_1192;
    _T_1194 <= _T_1193;
    _T_1195 <= _T_1194;
    _T_1196 <= _T_1195;
    _T_1197 <= _T_1196;
    _T_1198 <= _T_1197;
    _T_1199 <= _T_1198;
    _T_1200 <= _T_1199;
    _T_1201 <= _T_1200;
    _T_1202 <= _T_1201;
    _T_1203 <= _T_1202;
    _T_1204 <= _T_1203;
    _T_1205 <= _T_1204;
    _T_1206 <= _T_1205;
    _T_1207 <= _T_1206;
    _T_1208 <= _T_1207;
    _T_1209 <= _T_1208;
    _T_1210 <= _T_1209;
    _T_1211 <= _T_1210;
    _T_1212 <= _T_1211;
    _T_1213 <= _T_1212;
    _T_1214 <= _T_1213;
    _T_1215 <= _T_1214;
    _T_1216 <= _T_1215;
    _T_1217 <= _T_1216;
    _T_1218 <= _T_1217;
    _T_1219 <= _T_1218;
    _T_1220 <= _T_1219;
    _T_1221 <= _T_1220;
    _T_1222 <= _T_1221;
    _T_1223 <= _T_1222;
    _T_1224 <= _T_1223;
    _T_1225 <= _T_1224;
    _T_1226 <= _T_1225;
    _T_1227 <= _T_1226;
    _T_1228 <= _T_1227;
    _T_1229 <= _T_1228;
    _T_1230 <= _T_1229;
    _T_1231 <= _T_1230;
    _T_1232 <= _T_1231;
    _T_1233 <= _T_1232;
    _T_1234 <= _T_1233;
    _T_1235 <= _T_1234;
    _T_1236 <= _T_1235;
    _T_1237 <= _T_1236;
    _T_1238 <= _T_1237;
    _T_1239 <= _T_1238;
    _T_1240 <= _T_1239;
    _T_1241 <= _T_1240;
    _T_1242 <= _T_1241;
    _T_1243 <= _T_1242;
    _T_1244 <= _T_1243;
    _T_1245 <= _T_1244;
    _T_1246 <= _T_1245;
    _T_1247 <= _T_1246;
    _T_1248 <= _T_1247;
    _T_1249 <= _T_1248;
    _T_1250 <= _T_1249;
    _T_1251 <= _T_1250;
    _T_1252 <= _T_1251;
    _T_1253 <= _T_1252;
    _T_1254 <= _T_1253;
    _T_1255 <= _T_1254;
    _T_1256 <= _T_1255;
    _T_1257 <= _T_1256;
    _T_1258 <= _T_1257;
    _T_1259 <= _T_1258;
    _T_1260 <= _T_1259;
    _T_1261 <= _T_1260;
    _T_1262 <= _T_1261;
    _T_1263 <= _T_1262;
    _T_1264 <= _T_1263;
    _T_1265 <= _T_1264;
    _T_1266 <= _T_1265;
    _T_1267 <= _T_1266;
    _T_1268 <= _T_1267;
    _T_1269 <= _T_1268;
    _T_1270 <= _T_1269;
    _T_1271 <= _T_1270;
    _T_1272 <= _T_1271;
    _T_1273 <= _T_1272;
    _T_1274 <= _T_1273;
    _T_1275 <= _T_1274;
    _T_1276 <= _T_1275;
    _T_1277 <= _T_1276;
    _T_1278 <= _T_1277;
    _T_1279 <= _T_1278;
    _T_1280 <= _T_1279;
    _T_1281 <= _T_1280;
    _T_1282 <= _T_1281;
    _T_1283 <= _T_1282;
    _T_1284 <= _T_1283;
    _T_1285 <= _T_1284;
    _T_1286 <= _T_1285;
    _T_1287 <= _T_1286;
    _T_1288 <= _T_1287;
    _T_1289 <= _T_1288;
    _T_1290 <= _T_1289;
    _T_1291 <= _T_1290;
    _T_1292 <= _T_1291;
    _T_1293 <= _T_1292;
    _T_1294 <= _T_1293;
    _T_1295 <= _T_1294;
    _T_1296 <= _T_1295;
    _T_1297 <= _T_1296;
    _T_1298 <= _T_1297;
    _T_1299 <= _T_1298;
    _T_1300 <= _T_1299;
    _T_1301 <= _T_1300;
    _T_1302 <= _T_1301;
    _T_1303 <= _T_1302;
    _T_1304 <= _T_1303;
    _T_1305 <= _T_1304;
    _T_1306 <= _T_1305;
    _T_1307 <= _T_1306;
    _T_1308 <= _T_1307;
    _T_1309 <= _T_1308;
    _T_1310 <= _T_1309;
    _T_1311 <= _T_1310;
    _T_1312 <= _T_1311;
    _T_1313 <= _T_1312;
    _T_1314 <= _T_1313;
    _T_1315 <= _T_1314;
    _T_1316 <= _T_1315;
    _T_1317 <= _T_1316;
    _T_1318 <= _T_1317;
    _T_1319 <= _T_1318;
    _T_1320 <= _T_1319;
    _T_1321 <= _T_1320;
    _T_1322 <= _T_1321;
    _T_1323 <= _T_1322;
    _T_1324 <= _T_1323;
    _T_1325 <= _T_1324;
    _T_1326 <= _T_1325;
    _T_1327 <= _T_1326;
    _T_1328 <= _T_1327;
    _T_1329 <= _T_1328;
    _T_1330 <= _T_1329;
    _T_1331 <= _T_1330;
    _T_1332 <= _T_1331;
    _T_1333 <= _T_1332;
    _T_1334 <= _T_1333;
    _T_1335 <= _T_1334;
    _T_1336 <= _T_1335;
    _T_1337 <= _T_1336;
    _T_1338 <= _T_1337;
    _T_1339 <= _T_1338;
    _T_1340 <= _T_1339;
    _T_1341 <= _T_1340;
    _T_1342 <= _T_1341;
    _T_1343 <= _T_1342;
    _T_1344 <= _T_1343;
    _T_1345 <= _T_1344;
    _T_1346 <= _T_1345;
    _T_1347 <= _T_1346;
    _T_1348 <= _T_1347;
    _T_1349 <= _T_1348;
    _T_1350 <= _T_1349;
    _T_1351 <= _T_1350;
    _T_1352 <= _T_1351;
    _T_1353 <= _T_1352;
    _T_1354 <= _T_1353;
    _T_1355 <= _T_1354;
    _T_1356 <= _T_1355;
    _T_1357 <= _T_1356;
    _T_1358 <= _T_1357;
    _T_1359 <= _T_1358;
    _T_1360 <= _T_1359;
    _T_1361 <= _T_1360;
    _T_1362 <= _T_1361;
    _T_1363 <= _T_1362;
    _T_1364 <= _T_1363;
    _T_1365 <= _T_1364;
    _T_1366 <= _T_1365;
    _T_1367 <= _T_1366;
    _T_1368 <= _T_1367;
    _T_1369 <= _T_1368;
    _T_1370 <= _T_1369;
    _T_1371 <= _T_1370;
    _T_1372 <= _T_1371;
    _T_1373 <= _T_1372;
    _T_1374 <= _T_1373;
    _T_1375 <= _T_1374;
    _T_1376 <= _T_1375;
    _T_1377 <= _T_1376;
    _T_1378 <= _T_1377;
    _T_1379 <= _T_1378;
    _T_1380 <= _T_1379;
    _T_1381 <= _T_1380;
    _T_1382 <= _T_1381;
    _T_1383 <= _T_1382;
    _T_1384 <= _T_1383;
    _T_1385 <= _T_1384;
    _T_1386 <= _T_1385;
    _T_1387 <= _T_1386;
    _T_1388 <= _T_1387;
    _T_1389 <= _T_1388;
    _T_1390 <= _T_1389;
    _T_1391 <= _T_1390;
    _T_1392 <= _T_1391;
    _T_1393 <= _T_1392;
    _T_1394 <= _T_1393;
    _T_1395 <= _T_1394;
    _T_1396 <= _T_1395;
    _T_1397 <= _T_1396;
    _T_1398 <= _T_1397;
    _T_1399 <= _T_1398;
    _T_1400 <= _T_1399;
    _T_1401 <= _T_1400;
    _T_1402 <= _T_1401;
    _T_1403 <= _T_1402;
    _T_1404 <= _T_1403;
    _T_1405 <= _T_1404;
    _T_1406 <= _T_1405;
    _T_1407 <= _T_1406;
    _T_1408 <= _T_1407;
    _T_1409 <= _T_1408;
    _T_1410 <= _T_1409;
    _T_1411 <= _T_1410;
    _T_1412 <= _T_1411;
    _T_1413 <= _T_1412;
    _T_1414 <= _T_1413;
    _T_1415 <= _T_1414;
    _T_1416 <= _T_1415;
    _T_1417 <= _T_1416;
    _T_1418 <= _T_1417;
    _T_1419 <= _T_1418;
    _T_1420 <= _T_1419;
    _T_1421 <= _T_1420;
    _T_1422 <= _T_1421;
    _T_1423 <= _T_1422;
    _T_1424 <= _T_1423;
    _T_1425 <= _T_1424;
    _T_1426 <= _T_1425;
    _T_1427 <= _T_1426;
    _T_1428 <= _T_1427;
    _T_1429 <= _T_1428;
    _T_1430 <= _T_1429;
    _T_1431 <= _T_1430;
    _T_1432 <= _T_1431;
    _T_1433 <= _T_1432;
    _T_1434 <= _T_1433;
    _T_1435 <= _T_1434;
    _T_1436 <= _T_1435;
    _T_1437 <= _T_1436;
    _T_1438 <= _T_1437;
    _T_1439 <= _T_1438;
    _T_1440 <= _T_1439;
    _T_1441 <= _T_1440;
    _T_1442 <= _T_1441;
    _T_1443 <= _T_1442;
    _T_1444 <= _T_1443;
    _T_1445 <= _T_1444;
    _T_1446 <= _T_1445;
    _T_1447 <= _T_1446;
    _T_1448 <= _T_1447;
    _T_1449 <= _T_1448;
    _T_1450 <= _T_1449;
    _T_1451 <= _T_1450;
    _T_1452 <= _T_1451;
    _T_1453 <= _T_1452;
    _T_1454 <= _T_1453;
    _T_1455 <= _T_1454;
    _T_1456 <= _T_1455;
    _T_1457 <= _T_1456;
    _T_1458 <= _T_1457;
    _T_1459 <= _T_1458;
    _T_1460 <= _T_1459;
    _T_1461 <= _T_1460;
    _T_1462 <= _T_1461;
    _T_1463 <= _T_1462;
    _T_1464 <= _T_1463;
    _T_1465 <= _T_1464;
    _T_1466 <= _T_1465;
    _T_1467 <= _T_1466;
    _T_1468 <= _T_1467;
    _T_1469 <= _T_1468;
    _T_1470 <= _T_1469;
    _T_1471 <= _T_1470;
    _T_1472 <= _T_1471;
    _T_1473 <= _T_1472;
    _T_1474 <= _T_1473;
    _T_1475 <= _T_1474;
    _T_1476 <= _T_1475;
    _T_1477 <= _T_1476;
    _T_1478 <= _T_1477;
    _T_1479 <= _T_1478;
    _T_1480 <= _T_1479;
    _T_1481 <= _T_1480;
    _T_1482 <= _T_1481;
    _T_1483 <= _T_1482;
    _T_1484 <= _T_1483;
    _T_1485 <= _T_1484;
    _T_1486 <= _T_1485;
    _T_1487 <= _T_1486;
    _T_1488 <= _T_1487;
    _T_1489 <= _T_1488;
    _T_1490 <= _T_1489;
    _T_1491 <= _T_1490;
    _T_1492 <= _T_1491;
    _T_1493 <= _T_1492;
    _T_1494 <= _T_1493;
    _T_1495 <= _T_1494;
    _T_1496 <= _T_1495;
    _T_1497 <= _T_1496;
    _T_1498 <= _T_1497;
    _T_1499 <= io_din_valid;
    _T_1500 <= _T_1499;
    _T_1501 <= _T_1500;
    _T_1502 <= _T_1501;
    _T_1503 <= _T_1502;
    _T_1504 <= _T_1503;
    _T_1505 <= _T_1504;
    _T_1506 <= _T_1505;
    _T_1507 <= _T_1506;
    _T_1508 <= _T_1507;
    _T_1509 <= _T_1508;
    _T_1510 <= _T_1509;
    _T_1511 <= _T_1510;
    _T_1512 <= _T_1511;
    _T_1513 <= _T_1512;
    _T_1514 <= _T_1513;
    _T_1515 <= _T_1514;
    _T_1516 <= _T_1515;
    _T_1517 <= _T_1516;
    _T_1518 <= _T_1517;
    _T_1519 <= _T_1518;
    _T_1520 <= _T_1519;
    _T_1521 <= _T_1520;
    _T_1522 <= _T_1521;
    _T_1523 <= _T_1522;
    _T_1524 <= _T_1523;
    _T_1525 <= _T_1524;
    _T_1526 <= _T_1525;
    _T_1527 <= _T_1526;
    _T_1528 <= _T_1527;
    _T_1529 <= _T_1528;
    _T_1530 <= _T_1529;
    _T_1531 <= _T_1530;
    _T_1532 <= _T_1531;
    _T_1533 <= _T_1532;
    _T_1534 <= _T_1533;
    _T_1535 <= _T_1534;
    _T_1536 <= _T_1535;
    _T_1537 <= _T_1536;
    _T_1538 <= _T_1537;
    _T_1539 <= _T_1538;
    _T_1540 <= _T_1539;
    _T_1541 <= _T_1540;
    _T_1542 <= _T_1541;
    _T_1543 <= _T_1542;
    _T_1544 <= _T_1543;
    _T_1545 <= _T_1544;
    _T_1546 <= _T_1545;
    _T_1547 <= _T_1546;
    _T_1548 <= _T_1547;
    _T_1549 <= _T_1548;
    _T_1550 <= _T_1549;
    _T_1551 <= _T_1550;
    _T_1552 <= _T_1551;
    _T_1553 <= _T_1552;
    _T_1554 <= _T_1553;
    _T_1555 <= _T_1554;
    _T_1556 <= _T_1555;
    _T_1557 <= _T_1556;
    _T_1558 <= _T_1557;
    _T_1559 <= _T_1558;
    _T_1560 <= _T_1559;
    _T_1561 <= _T_1560;
    _T_1562 <= _T_1561;
    _T_1563 <= _T_1562;
    _T_1564 <= _T_1563;
    _T_1565 <= _T_1564;
    _T_1566 <= _T_1565;
    _T_1567 <= _T_1566;
    _T_1568 <= _T_1567;
    _T_1569 <= _T_1568;
    _T_1570 <= _T_1569;
    _T_1571 <= _T_1570;
    _T_1572 <= _T_1571;
    _T_1573 <= _T_1572;
    _T_1574 <= _T_1573;
    _T_1575 <= _T_1574;
    _T_1576 <= _T_1575;
    _T_1577 <= _T_1576;
    _T_1578 <= _T_1577;
    _T_1579 <= _T_1578;
    _T_1580 <= _T_1579;
    _T_1581 <= _T_1580;
    _T_1582 <= _T_1581;
    _T_1583 <= _T_1582;
    _T_1584 <= _T_1583;
    _T_1585 <= _T_1584;
    _T_1586 <= _T_1585;
    _T_1587 <= _T_1586;
    _T_1588 <= _T_1587;
    _T_1589 <= _T_1588;
    _T_1590 <= _T_1589;
    _T_1591 <= _T_1590;
    _T_1592 <= _T_1591;
    _T_1593 <= _T_1592;
    _T_1594 <= _T_1593;
    _T_1595 <= _T_1594;
    _T_1596 <= _T_1595;
    _T_1597 <= _T_1596;
    _T_1598 <= _T_1597;
    _T_1599 <= _T_1598;
    _T_1600 <= _T_1599;
    _T_1601 <= _T_1600;
    _T_1602 <= _T_1601;
    _T_1603 <= _T_1602;
    _T_1604 <= _T_1603;
    _T_1605 <= _T_1604;
    _T_1606 <= _T_1605;
    _T_1607 <= _T_1606;
    _T_1608 <= _T_1607;
    _T_1609 <= _T_1608;
    _T_1610 <= _T_1609;
    _T_1611 <= _T_1610;
    _T_1612 <= _T_1611;
    _T_1613 <= _T_1612;
    _T_1614 <= _T_1613;
    _T_1615 <= _T_1614;
    _T_1616 <= _T_1615;
    _T_1617 <= _T_1616;
    _T_1618 <= _T_1617;
    _T_1619 <= _T_1618;
    _T_1620 <= _T_1619;
    _T_1621 <= _T_1620;
    _T_1622 <= _T_1621;
    _T_1623 <= _T_1622;
    _T_1624 <= _T_1623;
    _T_1625 <= _T_1624;
    _T_1626 <= _T_1625;
    _T_1627 <= _T_1626;
    _T_1628 <= _T_1627;
    _T_1629 <= _T_1628;
    _T_1630 <= _T_1629;
    _T_1631 <= _T_1630;
    _T_1632 <= _T_1631;
    _T_1633 <= _T_1632;
    _T_1634 <= _T_1633;
    _T_1635 <= _T_1634;
    _T_1636 <= _T_1635;
    _T_1637 <= _T_1636;
    _T_1638 <= _T_1637;
    _T_1639 <= _T_1638;
    _T_1640 <= _T_1639;
    _T_1641 <= _T_1640;
    _T_1642 <= _T_1641;
    _T_1643 <= _T_1642;
    _T_1644 <= _T_1643;
    _T_1645 <= _T_1644;
    _T_1646 <= _T_1645;
    _T_1647 <= _T_1646;
    _T_1648 <= _T_1647;
    _T_1649 <= _T_1648;
    _T_1650 <= _T_1649;
    _T_1651 <= _T_1650;
    _T_1652 <= _T_1651;
    _T_1653 <= _T_1652;
    _T_1654 <= _T_1653;
    _T_1655 <= _T_1654;
    _T_1656 <= _T_1655;
    _T_1657 <= _T_1656;
    _T_1658 <= _T_1657;
    _T_1659 <= _T_1658;
    _T_1660 <= _T_1659;
    _T_1661 <= _T_1660;
    _T_1662 <= _T_1661;
    _T_1663 <= _T_1662;
    _T_1664 <= _T_1663;
    _T_1665 <= _T_1664;
    _T_1666 <= _T_1665;
    _T_1667 <= _T_1666;
    _T_1668 <= _T_1667;
    _T_1669 <= _T_1668;
    _T_1670 <= _T_1669;
    _T_1671 <= _T_1670;
    _T_1672 <= _T_1671;
    _T_1673 <= _T_1672;
    _T_1674 <= _T_1673;
    _T_1675 <= _T_1674;
    _T_1676 <= _T_1675;
    _T_1677 <= _T_1676;
    _T_1678 <= _T_1677;
    _T_1679 <= _T_1678;
    _T_1680 <= _T_1679;
    _T_1681 <= _T_1680;
    _T_1682 <= _T_1681;
    _T_1683 <= _T_1682;
    _T_1684 <= _T_1683;
    _T_1685 <= _T_1684;
    _T_1686 <= _T_1685;
    _T_1687 <= _T_1686;
    _T_1688 <= _T_1687;
    _T_1689 <= _T_1688;
    _T_1690 <= _T_1689;
    _T_1691 <= _T_1690;
    _T_1692 <= _T_1691;
    _T_1693 <= _T_1692;
    _T_1694 <= _T_1693;
    _T_1695 <= _T_1694;
    _T_1696 <= _T_1695;
    _T_1697 <= _T_1696;
    _T_1698 <= _T_1697;
    _T_1699 <= _T_1698;
    _T_1700 <= _T_1699;
    _T_1701 <= _T_1700;
    _T_1702 <= _T_1701;
    _T_1703 <= _T_1702;
    _T_1704 <= _T_1703;
    _T_1705 <= _T_1704;
    _T_1706 <= _T_1705;
    _T_1707 <= _T_1706;
    _T_1708 <= _T_1707;
    _T_1709 <= _T_1708;
    _T_1710 <= _T_1709;
    _T_1711 <= _T_1710;
    _T_1712 <= _T_1711;
    _T_1713 <= _T_1712;
    _T_1714 <= _T_1713;
    _T_1715 <= _T_1714;
    _T_1716 <= _T_1715;
    _T_1717 <= _T_1716;
    _T_1718 <= _T_1717;
    _T_1719 <= _T_1718;
    _T_1720 <= _T_1719;
    _T_1721 <= _T_1720;
    _T_1722 <= _T_1721;
    _T_1723 <= _T_1722;
    _T_1724 <= _T_1723;
    _T_1725 <= _T_1724;
    _T_1726 <= _T_1725;
    _T_1727 <= _T_1726;
    _T_1728 <= _T_1727;
    _T_1729 <= _T_1728;
    _T_1730 <= _T_1729;
    _T_1731 <= _T_1730;
    _T_1732 <= _T_1731;
    _T_1733 <= _T_1732;
    _T_1734 <= _T_1733;
    _T_1735 <= _T_1734;
    _T_1736 <= _T_1735;
    _T_1737 <= _T_1736;
    _T_1738 <= _T_1737;
    _T_1739 <= _T_1738;
    _T_1740 <= _T_1739;
    _T_1741 <= _T_1740;
    _T_1742 <= _T_1741;
    _T_1743 <= _T_1742;
    _T_1744 <= _T_1743;
    _T_1745 <= _T_1744;
    _T_1746 <= _T_1745;
    _T_1747 <= _T_1746;
    _T_1748 <= _T_1747;
    _T_1749 <= _T_1748;
    _T_1750 <= _T_1749;
    _T_1751 <= _T_1750;
    _T_1752 <= _T_1751;
    _T_1753 <= _T_1752;
    _T_1754 <= _T_1753;
    _T_1755 <= _T_1754;
    _T_1756 <= _T_1755;
    _T_1757 <= _T_1756;
    _T_1758 <= _T_1757;
    _T_1759 <= _T_1758;
    _T_1760 <= _T_1759;
    _T_1761 <= _T_1760;
    _T_1762 <= _T_1761;
    _T_1763 <= _T_1762;
    _T_1764 <= _T_1763;
    _T_1765 <= _T_1764;
    _T_1766 <= _T_1765;
    _T_1767 <= _T_1766;
    _T_1768 <= _T_1767;
    _T_1769 <= _T_1768;
    _T_1770 <= _T_1769;
    _T_1771 <= _T_1770;
    _T_1772 <= _T_1771;
    _T_1773 <= _T_1772;
    _T_1774 <= _T_1773;
    _T_1775 <= _T_1774;
    _T_1776 <= _T_1775;
    _T_1777 <= _T_1776;
    _T_1778 <= _T_1777;
    _T_1779 <= _T_1778;
    _T_1780 <= _T_1779;
    _T_1781 <= _T_1780;
    _T_1782 <= _T_1781;
    _T_1783 <= _T_1782;
    _T_1784 <= _T_1783;
    _T_1785 <= _T_1784;
    _T_1786 <= _T_1785;
    _T_1787 <= _T_1786;
    _T_1788 <= _T_1787;
    _T_1789 <= _T_1788;
    _T_1790 <= _T_1789;
    _T_1791 <= _T_1790;
    _T_1792 <= _T_1791;
    _T_1793 <= _T_1792;
    _T_1794 <= _T_1793;
    _T_1795 <= _T_1794;
    _T_1796 <= _T_1795;
    _T_1797 <= _T_1796;
    _T_1798 <= _T_1797;
    _T_1799 <= _T_1798;
    _T_1800 <= _T_1799;
    _T_1801 <= _T_1800;
    _T_1802 <= _T_1801;
    _T_1803 <= _T_1802;
    _T_1804 <= _T_1803;
    _T_1805 <= _T_1804;
    _T_1806 <= _T_1805;
    _T_1807 <= _T_1806;
    _T_1808 <= _T_1807;
    _T_1809 <= _T_1808;
    _T_1810 <= _T_1809;
    _T_1811 <= _T_1810;
    _T_1812 <= _T_1811;
    _T_1813 <= _T_1812;
    _T_1814 <= _T_1813;
    _T_1815 <= _T_1814;
    _T_1816 <= _T_1815;
    _T_1817 <= _T_1816;
    _T_1818 <= _T_1817;
    _T_1819 <= _T_1818;
    _T_1820 <= _T_1819;
    _T_1821 <= _T_1820;
    _T_1822 <= _T_1821;
    _T_1823 <= _T_1822;
    _T_1824 <= _T_1823;
    _T_1825 <= _T_1824;
    _T_1826 <= _T_1825;
    _T_1827 <= _T_1826;
    _T_1828 <= _T_1827;
    _T_1829 <= _T_1828;
    _T_1830 <= _T_1829;
    _T_1831 <= _T_1830;
    _T_1832 <= _T_1831;
    _T_1833 <= _T_1832;
    _T_1834 <= _T_1833;
    _T_1835 <= _T_1834;
    _T_1836 <= _T_1835;
    _T_1837 <= _T_1836;
    _T_1838 <= _T_1837;
    _T_1839 <= _T_1838;
    _T_1840 <= _T_1839;
    _T_1841 <= _T_1840;
    _T_1842 <= _T_1841;
    _T_1843 <= _T_1842;
    _T_1844 <= _T_1843;
    _T_1845 <= _T_1844;
    _T_1846 <= _T_1845;
    _T_1847 <= _T_1846;
    _T_1848 <= _T_1847;
    _T_1849 <= _T_1848;
    _T_1850 <= _T_1849;
    _T_1851 <= _T_1850;
    _T_1852 <= _T_1851;
    _T_1853 <= _T_1852;
    _T_1854 <= _T_1853;
    _T_1855 <= _T_1854;
    _T_1856 <= _T_1855;
    _T_1857 <= _T_1856;
    _T_1858 <= _T_1857;
    _T_1859 <= _T_1858;
    _T_1860 <= _T_1859;
    _T_1861 <= _T_1860;
    _T_1862 <= _T_1861;
    _T_1863 <= _T_1862;
    _T_1864 <= _T_1863;
    _T_1865 <= _T_1864;
    _T_1866 <= _T_1865;
    _T_1867 <= _T_1866;
    _T_1868 <= _T_1867;
    _T_1869 <= _T_1868;
    _T_1870 <= _T_1869;
    _T_1871 <= _T_1870;
    _T_1872 <= _T_1871;
    _T_1873 <= _T_1872;
    _T_1874 <= _T_1873;
    _T_1875 <= _T_1874;
    _T_1876 <= _T_1875;
    _T_1877 <= _T_1876;
    _T_1878 <= _T_1877;
    _T_1879 <= _T_1878;
    _T_1880 <= _T_1879;
    _T_1881 <= _T_1880;
    _T_1882 <= _T_1881;
    _T_1883 <= _T_1882;
    _T_1884 <= _T_1883;
    _T_1885 <= _T_1884;
    _T_1886 <= _T_1885;
    _T_1887 <= _T_1886;
    _T_1888 <= _T_1887;
    _T_1889 <= _T_1888;
    _T_1890 <= _T_1889;
    _T_1891 <= _T_1890;
    _T_1892 <= _T_1891;
    _T_1893 <= _T_1892;
    _T_1894 <= _T_1893;
    _T_1895 <= _T_1894;
    _T_1896 <= _T_1895;
    _T_1897 <= _T_1896;
    _T_1898 <= _T_1897;
    _T_1899 <= _T_1898;
    _T_1900 <= _T_1899;
    _T_1901 <= _T_1900;
    _T_1902 <= _T_1901;
    _T_1903 <= _T_1902;
    _T_1904 <= _T_1903;
    _T_1905 <= _T_1904;
    _T_1906 <= _T_1905;
    _T_1907 <= _T_1906;
    _T_1908 <= _T_1907;
    _T_1909 <= _T_1908;
    _T_1910 <= _T_1909;
    _T_1911 <= _T_1910;
    _T_1912 <= _T_1911;
    _T_1913 <= _T_1912;
    _T_1914 <= _T_1913;
    _T_1915 <= _T_1914;
    _T_1916 <= _T_1915;
    _T_1917 <= _T_1916;
    _T_1918 <= _T_1917;
    _T_1919 <= _T_1918;
    _T_1920 <= _T_1919;
    _T_1921 <= _T_1920;
    _T_1922 <= _T_1921;
    _T_1923 <= _T_1922;
    _T_1924 <= _T_1923;
    _T_1925 <= _T_1924;
    _T_1926 <= _T_1925;
    _T_1927 <= _T_1926;
    _T_1928 <= _T_1927;
    _T_1929 <= _T_1928;
    _T_1930 <= _T_1929;
    _T_1931 <= _T_1930;
    _T_1932 <= _T_1931;
    _T_1933 <= _T_1932;
    _T_1934 <= _T_1933;
    _T_1935 <= _T_1934;
    _T_1936 <= _T_1935;
    _T_1937 <= _T_1936;
    _T_1938 <= _T_1937;
    _T_1939 <= _T_1938;
    _T_1940 <= _T_1939;
    _T_1941 <= _T_1940;
    _T_1942 <= _T_1941;
    _T_1943 <= _T_1942;
    _T_1944 <= _T_1943;
    _T_1945 <= _T_1944;
    _T_1946 <= _T_1945;
    _T_1947 <= _T_1946;
    _T_1948 <= _T_1947;
    _T_1949 <= _T_1948;
    _T_1950 <= _T_1949;
    _T_1951 <= _T_1950;
    _T_1952 <= _T_1951;
    _T_1953 <= _T_1952;
    _T_1954 <= _T_1953;
    _T_1955 <= _T_1954;
    _T_1956 <= _T_1955;
    _T_1957 <= _T_1956;
    _T_1958 <= _T_1957;
    _T_1959 <= _T_1958;
    _T_1960 <= _T_1959;
    _T_1961 <= _T_1960;
    _T_1962 <= _T_1961;
    _T_1963 <= _T_1962;
    _T_1964 <= _T_1963;
    _T_1965 <= _T_1964;
    _T_1966 <= _T_1965;
    _T_1967 <= _T_1966;
    _T_1968 <= _T_1967;
    _T_1969 <= _T_1968;
    _T_1970 <= _T_1969;
    _T_1971 <= _T_1970;
    _T_1972 <= _T_1971;
    _T_1973 <= _T_1972;
    _T_1974 <= _T_1973;
    _T_1975 <= _T_1974;
    _T_1976 <= _T_1975;
    _T_1977 <= _T_1976;
    _T_1978 <= _T_1977;
    _T_1979 <= _T_1978;
    _T_1980 <= _T_1979;
    _T_1981 <= _T_1980;
    _T_1982 <= _T_1981;
    _T_1983 <= _T_1982;
    _T_1984 <= _T_1983;
    _T_1985 <= _T_1984;
    _T_1986 <= _T_1985;
    _T_1987 <= _T_1986;
    _T_1988 <= _T_1987;
    _T_1989 <= _T_1988;
    _T_1990 <= _T_1989;
    _T_1991 <= _T_1990;
    _T_1992 <= _T_1991;
    _T_1993 <= _T_1992;
    _T_1994 <= _T_1993;
    _T_1995 <= _T_1994;
    _T_1996 <= _T_1995;
    _T_1997 <= _T_1996;
    _T_1998 <= _T_1997;
    _T_1999 <= _T_1998;
    _T_2000 <= _T_1999;
    _T_2001 <= _T_2000;
    _T_2002 <= _T_2001;
    _T_2003 <= _T_2002;
    _T_2004 <= _T_2003;
    _T_2005 <= _T_2004;
    _T_2006 <= _T_2005;
    _T_2007 <= _T_2006;
    _T_2008 <= _T_2007;
    _T_2009 <= _T_2008;
    _T_2010 <= _T_2009;
    _T_2011 <= _T_2010;
    _T_2012 <= _T_2011;
    _T_2013 <= _T_2012;
    _T_2014 <= _T_2013;
    _T_2015 <= _T_2014;
    _T_2016 <= _T_2015;
    _T_2017 <= _T_2016;
    _T_2018 <= _T_2017;
    _T_2019 <= _T_2018;
    _T_2020 <= _T_2019;
    _T_2021 <= _T_2020;
    _T_2022 <= _T_2021;
    _T_2023 <= _T_2022;
    _T_2024 <= _T_2023;
    _T_2025 <= _T_2024;
    _T_2026 <= _T_2025;
    _T_2027 <= _T_2026;
    _T_2028 <= _T_2027;
    _T_2029 <= _T_2028;
    _T_2030 <= _T_2029;
    _T_2031 <= _T_2030;
    _T_2032 <= _T_2031;
    _T_2033 <= _T_2032;
    _T_2034 <= _T_2033;
    _T_2035 <= _T_2034;
    _T_2036 <= _T_2035;
    _T_2037 <= _T_2036;
    _T_2038 <= _T_2037;
    _T_2039 <= _T_2038;
    _T_2040 <= _T_2039;
    _T_2041 <= _T_2040;
    _T_2042 <= _T_2041;
    _T_2043 <= _T_2042;
    _T_2044 <= _T_2043;
    _T_2045 <= _T_2044;
    _T_2046 <= _T_2045;
    _T_2047 <= _T_2046;
    _T_2048 <= _T_2047;
    _T_2049 <= _T_2048;
    _T_2050 <= _T_2049;
    _T_2051 <= _T_2050;
    _T_2052 <= _T_2051;
    _T_2053 <= _T_2052;
    _T_2054 <= _T_2053;
    _T_2055 <= _T_2054;
    _T_2056 <= _T_2055;
    _T_2057 <= _T_2056;
    _T_2058 <= _T_2057;
    _T_2059 <= _T_2058;
    _T_2060 <= _T_2059;
    _T_2061 <= _T_2060;
    _T_2062 <= _T_2061;
    _T_2063 <= _T_2062;
    _T_2064 <= _T_2063;
    _T_2065 <= _T_2064;
    _T_2066 <= _T_2065;
    _T_2067 <= _T_2066;
    _T_2068 <= _T_2067;
    _T_2069 <= _T_2068;
    _T_2070 <= _T_2069;
    _T_2071 <= _T_2070;
    _T_2072 <= _T_2071;
    _T_2073 <= _T_2072;
    _T_2074 <= _T_2073;
    _T_2075 <= _T_2074;
    _T_2076 <= _T_2075;
    _T_2077 <= _T_2076;
    _T_2078 <= _T_2077;
    _T_2079 <= _T_2078;
    _T_2080 <= _T_2079;
    _T_2081 <= _T_2080;
    _T_2082 <= _T_2081;
    _T_2083 <= _T_2082;
    _T_2084 <= _T_2083;
    _T_2085 <= _T_2084;
    _T_2086 <= _T_2085;
    _T_2087 <= _T_2086;
    _T_2088 <= _T_2087;
    _T_2089 <= _T_2088;
    _T_2090 <= _T_2089;
    _T_2091 <= _T_2090;
    _T_2092 <= _T_2091;
    _T_2093 <= _T_2092;
    _T_2094 <= _T_2093;
    _T_2095 <= _T_2094;
    _T_2096 <= _T_2095;
    _T_2097 <= _T_2096;
    _T_2098 <= _T_2097;
    _T_2099 <= _T_2098;
    _T_2100 <= _T_2099;
    _T_2101 <= _T_2100;
    _T_2102 <= _T_2101;
    _T_2103 <= _T_2102;
    _T_2104 <= _T_2103;
    _T_2105 <= _T_2104;
    _T_2106 <= _T_2105;
    _T_2107 <= _T_2106;
    _T_2108 <= _T_2107;
    _T_2109 <= _T_2108;
    _T_2110 <= _T_2109;
    _T_2111 <= _T_2110;
    _T_2112 <= _T_2111;
    _T_2113 <= _T_2112;
    _T_2114 <= _T_2113;
    _T_2115 <= _T_2114;
    _T_2116 <= _T_2115;
    _T_2117 <= _T_2116;
    _T_2118 <= _T_2117;
    _T_2119 <= _T_2118;
    _T_2120 <= _T_2119;
    _T_2121 <= _T_2120;
    _T_2122 <= _T_2121;
    _T_2123 <= _T_2122;
    _T_2124 <= _T_2123;
    _T_2125 <= _T_2124;
    _T_2126 <= _T_2125;
    _T_2127 <= _T_2126;
    _T_2128 <= _T_2127;
    _T_2129 <= _T_2128;
    _T_2130 <= _T_2129;
    _T_2131 <= _T_2130;
    _T_2132 <= _T_2131;
    _T_2133 <= _T_2132;
    _T_2134 <= _T_2133;
    _T_2135 <= _T_2134;
    _T_2136 <= _T_2135;
    _T_2137 <= _T_2136;
    _T_2138 <= _T_2137;
    _T_2139 <= _T_2138;
    _T_2140 <= _T_2139;
    _T_2141 <= _T_2140;
    _T_2142 <= _T_2141;
    _T_2143 <= _T_2142;
    _T_2144 <= _T_2143;
    _T_2145 <= _T_2144;
    _T_2146 <= _T_2145;
    _T_2147 <= _T_2146;
    _T_2148 <= _T_2147;
    _T_2149 <= _T_2148;
    _T_2150 <= _T_2149;
    _T_2151 <= _T_2150;
    _T_2152 <= _T_2151;
    _T_2153 <= _T_2152;
    _T_2154 <= _T_2153;
    _T_2155 <= _T_2154;
    _T_2156 <= _T_2155;
    _T_2157 <= _T_2156;
    _T_2158 <= _T_2157;
    _T_2159 <= _T_2158;
    _T_2160 <= _T_2159;
    _T_2161 <= _T_2160;
    _T_2162 <= _T_2161;
    _T_2163 <= _T_2162;
    _T_2164 <= _T_2163;
    _T_2165 <= _T_2164;
    _T_2166 <= _T_2165;
    _T_2167 <= _T_2166;
    _T_2168 <= _T_2167;
    _T_2169 <= _T_2168;
    _T_2170 <= _T_2169;
    _T_2171 <= _T_2170;
    _T_2172 <= _T_2171;
    _T_2173 <= _T_2172;
    _T_2174 <= _T_2173;
    _T_2175 <= _T_2174;
    _T_2176 <= _T_2175;
    _T_2177 <= _T_2176;
    _T_2178 <= _T_2177;
    _T_2179 <= _T_2178;
    _T_2180 <= _T_2179;
    _T_2181 <= _T_2180;
    _T_2182 <= _T_2181;
    _T_2183 <= _T_2182;
    _T_2184 <= _T_2183;
    _T_2185 <= _T_2184;
    _T_2186 <= _T_2185;
    _T_2187 <= _T_2186;
    _T_2188 <= _T_2187;
    _T_2189 <= _T_2188;
    _T_2190 <= _T_2189;
    _T_2191 <= _T_2190;
    _T_2192 <= _T_2191;
    _T_2193 <= _T_2192;
    _T_2194 <= _T_2193;
    _T_2195 <= _T_2194;
    _T_2196 <= _T_2195;
    _T_2197 <= _T_2196;
    _T_2198 <= _T_2197;
    _T_2199 <= _T_2198;
    _T_2200 <= _T_2199;
    _T_2201 <= _T_2200;
    _T_2202 <= _T_2201;
    _T_2203 <= _T_2202;
    _T_2204 <= _T_2203;
    _T_2205 <= _T_2204;
    _T_2206 <= _T_2205;
    _T_2207 <= _T_2206;
    _T_2208 <= _T_2207;
    _T_2209 <= _T_2208;
    _T_2210 <= _T_2209;
    _T_2211 <= _T_2210;
    _T_2212 <= _T_2211;
    _T_2213 <= _T_2212;
    _T_2214 <= _T_2213;
    _T_2215 <= _T_2214;
    _T_2216 <= _T_2215;
    _T_2217 <= _T_2216;
    _T_2218 <= _T_2217;
    _T_2219 <= _T_2218;
    _T_2220 <= _T_2219;
    _T_2221 <= _T_2220;
    _T_2222 <= _T_2221;
    _T_2223 <= _T_2222;
    _T_2224 <= _T_2223;
    _T_2225 <= _T_2224;
    _T_2226 <= _T_2225;
    _T_2227 <= _T_2226;
    _T_2228 <= _T_2227;
    _T_2229 <= _T_2228;
    _T_2230 <= _T_2229;
    _T_2231 <= _T_2230;
    _T_2232 <= _T_2231;
    _T_2233 <= _T_2232;
    _T_2234 <= _T_2233;
    _T_2235 <= _T_2234;
    _T_2236 <= _T_2235;
    _T_2237 <= _T_2236;
    _T_2238 <= _T_2237;
    _T_2239 <= _T_2238;
    _T_2240 <= _T_2239;
    _T_2241 <= _T_2240;
    _T_2242 <= _T_2241;
    _T_2243 <= _T_2242;
    _T_2244 <= _T_2243;
    _T_2245 <= _T_2244;
    _T_2246 <= _T_2245;
    _T_2247 <= _T_2246;
    _T_2248 <= _T_2247;
    _T_2249 <= _T_2248;
    _T_2250 <= _T_2249;
    _T_2251 <= _T_2250;
    _T_2252 <= _T_2251;
    _T_2253 <= _T_2252;
    _T_2254 <= _T_2253;
    _T_2255 <= _T_2254;
    _T_2256 <= _T_2255;
    _T_2257 <= _T_2256;
    _T_2258 <= _T_2257;
    _T_2259 <= _T_2258;
    _T_2260 <= _T_2259;
    _T_2261 <= _T_2260;
    _T_2262 <= _T_2261;
    _T_2263 <= _T_2262;
    _T_2264 <= _T_2263;
    _T_2265 <= _T_2264;
    _T_2266 <= _T_2265;
  end
endmodule
module Reorder(
  input         clock,
  input         reset,
  input  [31:0] io_in1_re,
  input  [31:0] io_in1_im,
  input  [31:0] io_in2_re,
  input  [31:0] io_in2_im,
  input         io_in_valid,
  output [31:0] io_out_re,
  output [31:0] io_out_im,
  output        io_out_valid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] rambank0_re [0:255]; // @[Reorder.scala 20:21]
  wire [31:0] rambank0_re__T_845_data; // @[Reorder.scala 20:21]
  wire [7:0] rambank0_re__T_845_addr; // @[Reorder.scala 20:21]
  wire [31:0] rambank0_re__T_69_data; // @[Reorder.scala 20:21]
  wire [7:0] rambank0_re__T_69_addr; // @[Reorder.scala 20:21]
  wire  rambank0_re__T_69_mask; // @[Reorder.scala 20:21]
  wire  rambank0_re__T_69_en; // @[Reorder.scala 20:21]
  reg [31:0] rambank0_im [0:255]; // @[Reorder.scala 20:21]
  wire [31:0] rambank0_im__T_845_data; // @[Reorder.scala 20:21]
  wire [7:0] rambank0_im__T_845_addr; // @[Reorder.scala 20:21]
  wire [31:0] rambank0_im__T_69_data; // @[Reorder.scala 20:21]
  wire [7:0] rambank0_im__T_69_addr; // @[Reorder.scala 20:21]
  wire  rambank0_im__T_69_mask; // @[Reorder.scala 20:21]
  wire  rambank0_im__T_69_en; // @[Reorder.scala 20:21]
  reg [31:0] rambank1_re [0:255]; // @[Reorder.scala 21:21]
  wire [31:0] rambank1_re__T_847_data; // @[Reorder.scala 21:21]
  wire [7:0] rambank1_re__T_847_addr; // @[Reorder.scala 21:21]
  wire [31:0] rambank1_re__T_71_data; // @[Reorder.scala 21:21]
  wire [7:0] rambank1_re__T_71_addr; // @[Reorder.scala 21:21]
  wire  rambank1_re__T_71_mask; // @[Reorder.scala 21:21]
  wire  rambank1_re__T_71_en; // @[Reorder.scala 21:21]
  reg [31:0] rambank1_im [0:255]; // @[Reorder.scala 21:21]
  wire [31:0] rambank1_im__T_847_data; // @[Reorder.scala 21:21]
  wire [7:0] rambank1_im__T_847_addr; // @[Reorder.scala 21:21]
  wire [31:0] rambank1_im__T_71_data; // @[Reorder.scala 21:21]
  wire [7:0] rambank1_im__T_71_addr; // @[Reorder.scala 21:21]
  wire  rambank1_im__T_71_mask; // @[Reorder.scala 21:21]
  wire  rambank1_im__T_71_en; // @[Reorder.scala 21:21]
  reg [7:0] in_counter; // @[Reorder.scala 25:27]
  reg [8:0] out_counter; // @[Reorder.scala 26:28]
  wire [8:0] _T = {in_counter,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_5 = {{4'd0}, _T[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_7 = {_T[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_9 = _T_7 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_10 = _T_5 | _T_9; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_787 = {{2'd0}, _T_10[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_15 = _GEN_787 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_17 = {_T_10[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_19 = _T_17 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_20 = _T_15 | _T_19; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_788 = {{1'd0}, _T_20[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_25 = _GEN_788 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_27 = {_T_20[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_29 = _T_27 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_30 = _T_25 | _T_29; // @[Bitwise.scala 103:39]
  wire [8:0] index1 = {_T_30,_T[8]}; // @[Cat.scala 29:58]
  wire [8:0] _T_32 = {in_counter,1'h1}; // @[Cat.scala 29:58]
  wire [7:0] _T_37 = {{4'd0}, _T_32[7:4]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_39 = {_T_32[3:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_41 = _T_39 & 8'hf0; // @[Bitwise.scala 103:75]
  wire [7:0] _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_789 = {{2'd0}, _T_42[7:2]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_47 = _GEN_789 & 8'h33; // @[Bitwise.scala 103:31]
  wire [7:0] _T_49 = {_T_42[5:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_51 = _T_49 & 8'hcc; // @[Bitwise.scala 103:75]
  wire [7:0] _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  wire [7:0] _GEN_790 = {{1'd0}, _T_52[7:1]}; // @[Bitwise.scala 103:31]
  wire [7:0] _T_57 = _GEN_790 & 8'h55; // @[Bitwise.scala 103:31]
  wire [7:0] _T_59 = {_T_52[6:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [7:0] _T_61 = _T_59 & 8'haa; // @[Bitwise.scala 103:75]
  wire [7:0] _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39]
  wire [8:0] index2 = {_T_62,_T_32[8]}; // @[Cat.scala 29:58]
  wire  _T_64 = ~io_out_valid; // @[Reorder.scala 29:23]
  wire  _T_65 = io_in_valid & _T_64; // @[Reorder.scala 29:20]
  wire [7:0] _T_67 = in_counter + 8'h1; // @[Reorder.scala 30:30]
  reg  _T_72; // @[Reg.scala 15:16]
  reg  _T_73; // @[Reg.scala 15:16]
  reg  _T_74; // @[Reg.scala 15:16]
  reg  _T_75; // @[Reg.scala 15:16]
  reg  _T_76; // @[Reg.scala 15:16]
  reg  _T_77; // @[Reg.scala 15:16]
  reg  _T_78; // @[Reg.scala 15:16]
  reg  _T_79; // @[Reg.scala 15:16]
  reg  _T_80; // @[Reg.scala 15:16]
  reg  _T_81; // @[Reg.scala 15:16]
  reg  _T_82; // @[Reg.scala 15:16]
  reg  _T_83; // @[Reg.scala 15:16]
  reg  _T_84; // @[Reg.scala 15:16]
  reg  _T_85; // @[Reg.scala 15:16]
  reg  _T_86; // @[Reg.scala 15:16]
  reg  _T_87; // @[Reg.scala 15:16]
  reg  _T_88; // @[Reg.scala 15:16]
  reg  _T_89; // @[Reg.scala 15:16]
  reg  _T_90; // @[Reg.scala 15:16]
  reg  _T_91; // @[Reg.scala 15:16]
  reg  _T_92; // @[Reg.scala 15:16]
  reg  _T_93; // @[Reg.scala 15:16]
  reg  _T_94; // @[Reg.scala 15:16]
  reg  _T_95; // @[Reg.scala 15:16]
  reg  _T_96; // @[Reg.scala 15:16]
  reg  _T_97; // @[Reg.scala 15:16]
  reg  _T_98; // @[Reg.scala 15:16]
  reg  _T_99; // @[Reg.scala 15:16]
  reg  _T_100; // @[Reg.scala 15:16]
  reg  _T_101; // @[Reg.scala 15:16]
  reg  _T_102; // @[Reg.scala 15:16]
  reg  _T_103; // @[Reg.scala 15:16]
  reg  _T_104; // @[Reg.scala 15:16]
  reg  _T_105; // @[Reg.scala 15:16]
  reg  _T_106; // @[Reg.scala 15:16]
  reg  _T_107; // @[Reg.scala 15:16]
  reg  _T_108; // @[Reg.scala 15:16]
  reg  _T_109; // @[Reg.scala 15:16]
  reg  _T_110; // @[Reg.scala 15:16]
  reg  _T_111; // @[Reg.scala 15:16]
  reg  _T_112; // @[Reg.scala 15:16]
  reg  _T_113; // @[Reg.scala 15:16]
  reg  _T_114; // @[Reg.scala 15:16]
  reg  _T_115; // @[Reg.scala 15:16]
  reg  _T_116; // @[Reg.scala 15:16]
  reg  _T_117; // @[Reg.scala 15:16]
  reg  _T_118; // @[Reg.scala 15:16]
  reg  _T_119; // @[Reg.scala 15:16]
  reg  _T_120; // @[Reg.scala 15:16]
  reg  _T_121; // @[Reg.scala 15:16]
  reg  _T_122; // @[Reg.scala 15:16]
  reg  _T_123; // @[Reg.scala 15:16]
  reg  _T_124; // @[Reg.scala 15:16]
  reg  _T_125; // @[Reg.scala 15:16]
  reg  _T_126; // @[Reg.scala 15:16]
  reg  _T_127; // @[Reg.scala 15:16]
  reg  _T_128; // @[Reg.scala 15:16]
  reg  _T_129; // @[Reg.scala 15:16]
  reg  _T_130; // @[Reg.scala 15:16]
  reg  _T_131; // @[Reg.scala 15:16]
  reg  _T_132; // @[Reg.scala 15:16]
  reg  _T_133; // @[Reg.scala 15:16]
  reg  _T_134; // @[Reg.scala 15:16]
  reg  _T_135; // @[Reg.scala 15:16]
  reg  _T_136; // @[Reg.scala 15:16]
  reg  _T_137; // @[Reg.scala 15:16]
  reg  _T_138; // @[Reg.scala 15:16]
  reg  _T_139; // @[Reg.scala 15:16]
  reg  _T_140; // @[Reg.scala 15:16]
  reg  _T_141; // @[Reg.scala 15:16]
  reg  _T_142; // @[Reg.scala 15:16]
  reg  _T_143; // @[Reg.scala 15:16]
  reg  _T_144; // @[Reg.scala 15:16]
  reg  _T_145; // @[Reg.scala 15:16]
  reg  _T_146; // @[Reg.scala 15:16]
  reg  _T_147; // @[Reg.scala 15:16]
  reg  _T_148; // @[Reg.scala 15:16]
  reg  _T_149; // @[Reg.scala 15:16]
  reg  _T_150; // @[Reg.scala 15:16]
  reg  _T_151; // @[Reg.scala 15:16]
  reg  _T_152; // @[Reg.scala 15:16]
  reg  _T_153; // @[Reg.scala 15:16]
  reg  _T_154; // @[Reg.scala 15:16]
  reg  _T_155; // @[Reg.scala 15:16]
  reg  _T_156; // @[Reg.scala 15:16]
  reg  _T_157; // @[Reg.scala 15:16]
  reg  _T_158; // @[Reg.scala 15:16]
  reg  _T_159; // @[Reg.scala 15:16]
  reg  _T_160; // @[Reg.scala 15:16]
  reg  _T_161; // @[Reg.scala 15:16]
  reg  _T_162; // @[Reg.scala 15:16]
  reg  _T_163; // @[Reg.scala 15:16]
  reg  _T_164; // @[Reg.scala 15:16]
  reg  _T_165; // @[Reg.scala 15:16]
  reg  _T_166; // @[Reg.scala 15:16]
  reg  _T_167; // @[Reg.scala 15:16]
  reg  _T_168; // @[Reg.scala 15:16]
  reg  _T_169; // @[Reg.scala 15:16]
  reg  _T_170; // @[Reg.scala 15:16]
  reg  _T_171; // @[Reg.scala 15:16]
  reg  _T_172; // @[Reg.scala 15:16]
  reg  _T_173; // @[Reg.scala 15:16]
  reg  _T_174; // @[Reg.scala 15:16]
  reg  _T_175; // @[Reg.scala 15:16]
  reg  _T_176; // @[Reg.scala 15:16]
  reg  _T_177; // @[Reg.scala 15:16]
  reg  _T_178; // @[Reg.scala 15:16]
  reg  _T_179; // @[Reg.scala 15:16]
  reg  _T_180; // @[Reg.scala 15:16]
  reg  _T_181; // @[Reg.scala 15:16]
  reg  _T_182; // @[Reg.scala 15:16]
  reg  _T_183; // @[Reg.scala 15:16]
  reg  _T_184; // @[Reg.scala 15:16]
  reg  _T_185; // @[Reg.scala 15:16]
  reg  _T_186; // @[Reg.scala 15:16]
  reg  _T_187; // @[Reg.scala 15:16]
  reg  _T_188; // @[Reg.scala 15:16]
  reg  _T_189; // @[Reg.scala 15:16]
  reg  _T_190; // @[Reg.scala 15:16]
  reg  _T_191; // @[Reg.scala 15:16]
  reg  _T_192; // @[Reg.scala 15:16]
  reg  _T_193; // @[Reg.scala 15:16]
  reg  _T_194; // @[Reg.scala 15:16]
  reg  _T_195; // @[Reg.scala 15:16]
  reg  _T_196; // @[Reg.scala 15:16]
  reg  _T_197; // @[Reg.scala 15:16]
  reg  _T_198; // @[Reg.scala 15:16]
  reg  _T_199; // @[Reg.scala 15:16]
  reg  _T_200; // @[Reg.scala 15:16]
  reg  _T_201; // @[Reg.scala 15:16]
  reg  _T_202; // @[Reg.scala 15:16]
  reg  _T_203; // @[Reg.scala 15:16]
  reg  _T_204; // @[Reg.scala 15:16]
  reg  _T_205; // @[Reg.scala 15:16]
  reg  _T_206; // @[Reg.scala 15:16]
  reg  _T_207; // @[Reg.scala 15:16]
  reg  _T_208; // @[Reg.scala 15:16]
  reg  _T_209; // @[Reg.scala 15:16]
  reg  _T_210; // @[Reg.scala 15:16]
  reg  _T_211; // @[Reg.scala 15:16]
  reg  _T_212; // @[Reg.scala 15:16]
  reg  _T_213; // @[Reg.scala 15:16]
  reg  _T_214; // @[Reg.scala 15:16]
  reg  _T_215; // @[Reg.scala 15:16]
  reg  _T_216; // @[Reg.scala 15:16]
  reg  _T_217; // @[Reg.scala 15:16]
  reg  _T_218; // @[Reg.scala 15:16]
  reg  _T_219; // @[Reg.scala 15:16]
  reg  _T_220; // @[Reg.scala 15:16]
  reg  _T_221; // @[Reg.scala 15:16]
  reg  _T_222; // @[Reg.scala 15:16]
  reg  _T_223; // @[Reg.scala 15:16]
  reg  _T_224; // @[Reg.scala 15:16]
  reg  _T_225; // @[Reg.scala 15:16]
  reg  _T_226; // @[Reg.scala 15:16]
  reg  _T_227; // @[Reg.scala 15:16]
  reg  _T_228; // @[Reg.scala 15:16]
  reg  _T_229; // @[Reg.scala 15:16]
  reg  _T_230; // @[Reg.scala 15:16]
  reg  _T_231; // @[Reg.scala 15:16]
  reg  _T_232; // @[Reg.scala 15:16]
  reg  _T_233; // @[Reg.scala 15:16]
  reg  _T_234; // @[Reg.scala 15:16]
  reg  _T_235; // @[Reg.scala 15:16]
  reg  _T_236; // @[Reg.scala 15:16]
  reg  _T_237; // @[Reg.scala 15:16]
  reg  _T_238; // @[Reg.scala 15:16]
  reg  _T_239; // @[Reg.scala 15:16]
  reg  _T_240; // @[Reg.scala 15:16]
  reg  _T_241; // @[Reg.scala 15:16]
  reg  _T_242; // @[Reg.scala 15:16]
  reg  _T_243; // @[Reg.scala 15:16]
  reg  _T_244; // @[Reg.scala 15:16]
  reg  _T_245; // @[Reg.scala 15:16]
  reg  _T_246; // @[Reg.scala 15:16]
  reg  _T_247; // @[Reg.scala 15:16]
  reg  _T_248; // @[Reg.scala 15:16]
  reg  _T_249; // @[Reg.scala 15:16]
  reg  _T_250; // @[Reg.scala 15:16]
  reg  _T_251; // @[Reg.scala 15:16]
  reg  _T_252; // @[Reg.scala 15:16]
  reg  _T_253; // @[Reg.scala 15:16]
  reg  _T_254; // @[Reg.scala 15:16]
  reg  _T_255; // @[Reg.scala 15:16]
  reg  _T_256; // @[Reg.scala 15:16]
  reg  _T_257; // @[Reg.scala 15:16]
  reg  _T_258; // @[Reg.scala 15:16]
  reg  _T_259; // @[Reg.scala 15:16]
  reg  _T_260; // @[Reg.scala 15:16]
  reg  _T_261; // @[Reg.scala 15:16]
  reg  _T_262; // @[Reg.scala 15:16]
  reg  _T_263; // @[Reg.scala 15:16]
  reg  _T_264; // @[Reg.scala 15:16]
  reg  _T_265; // @[Reg.scala 15:16]
  reg  _T_266; // @[Reg.scala 15:16]
  reg  _T_267; // @[Reg.scala 15:16]
  reg  _T_268; // @[Reg.scala 15:16]
  reg  _T_269; // @[Reg.scala 15:16]
  reg  _T_270; // @[Reg.scala 15:16]
  reg  _T_271; // @[Reg.scala 15:16]
  reg  _T_272; // @[Reg.scala 15:16]
  reg  _T_273; // @[Reg.scala 15:16]
  reg  _T_274; // @[Reg.scala 15:16]
  reg  _T_275; // @[Reg.scala 15:16]
  reg  _T_276; // @[Reg.scala 15:16]
  reg  _T_277; // @[Reg.scala 15:16]
  reg  _T_278; // @[Reg.scala 15:16]
  reg  _T_279; // @[Reg.scala 15:16]
  reg  _T_280; // @[Reg.scala 15:16]
  reg  _T_281; // @[Reg.scala 15:16]
  reg  _T_282; // @[Reg.scala 15:16]
  reg  _T_283; // @[Reg.scala 15:16]
  reg  _T_284; // @[Reg.scala 15:16]
  reg  _T_285; // @[Reg.scala 15:16]
  reg  _T_286; // @[Reg.scala 15:16]
  reg  _T_287; // @[Reg.scala 15:16]
  reg  _T_288; // @[Reg.scala 15:16]
  reg  _T_289; // @[Reg.scala 15:16]
  reg  _T_290; // @[Reg.scala 15:16]
  reg  _T_291; // @[Reg.scala 15:16]
  reg  _T_292; // @[Reg.scala 15:16]
  reg  _T_293; // @[Reg.scala 15:16]
  reg  _T_294; // @[Reg.scala 15:16]
  reg  _T_295; // @[Reg.scala 15:16]
  reg  _T_296; // @[Reg.scala 15:16]
  reg  _T_297; // @[Reg.scala 15:16]
  reg  _T_298; // @[Reg.scala 15:16]
  reg  _T_299; // @[Reg.scala 15:16]
  reg  _T_300; // @[Reg.scala 15:16]
  reg  _T_301; // @[Reg.scala 15:16]
  reg  _T_302; // @[Reg.scala 15:16]
  reg  _T_303; // @[Reg.scala 15:16]
  reg  _T_304; // @[Reg.scala 15:16]
  reg  _T_305; // @[Reg.scala 15:16]
  reg  _T_306; // @[Reg.scala 15:16]
  reg  _T_307; // @[Reg.scala 15:16]
  reg  _T_308; // @[Reg.scala 15:16]
  reg  _T_309; // @[Reg.scala 15:16]
  reg  _T_310; // @[Reg.scala 15:16]
  reg  _T_311; // @[Reg.scala 15:16]
  reg  _T_312; // @[Reg.scala 15:16]
  reg  _T_313; // @[Reg.scala 15:16]
  reg  _T_314; // @[Reg.scala 15:16]
  reg  _T_315; // @[Reg.scala 15:16]
  reg  _T_316; // @[Reg.scala 15:16]
  reg  _T_317; // @[Reg.scala 15:16]
  reg  _T_318; // @[Reg.scala 15:16]
  reg  _T_319; // @[Reg.scala 15:16]
  reg  _T_320; // @[Reg.scala 15:16]
  reg  _T_321; // @[Reg.scala 15:16]
  reg  _T_322; // @[Reg.scala 15:16]
  reg  _T_323; // @[Reg.scala 15:16]
  reg  _T_324; // @[Reg.scala 15:16]
  reg  _T_325; // @[Reg.scala 15:16]
  reg  _T_326; // @[Reg.scala 15:16]
  reg  _T_327; // @[Reg.scala 15:16]
  reg  _T_328; // @[Reg.scala 15:16]
  reg  _T_329; // @[Reg.scala 15:16]
  reg  _T_330; // @[Reg.scala 15:16]
  reg  _T_331; // @[Reg.scala 15:16]
  reg  _T_332; // @[Reg.scala 15:16]
  reg  _T_333; // @[Reg.scala 15:16]
  reg  _T_334; // @[Reg.scala 15:16]
  reg  _T_335; // @[Reg.scala 15:16]
  reg  _T_336; // @[Reg.scala 15:16]
  reg  _T_337; // @[Reg.scala 15:16]
  reg  _T_338; // @[Reg.scala 15:16]
  reg  _T_339; // @[Reg.scala 15:16]
  reg  _T_340; // @[Reg.scala 15:16]
  reg  _T_341; // @[Reg.scala 15:16]
  reg  _T_342; // @[Reg.scala 15:16]
  reg  _T_343; // @[Reg.scala 15:16]
  reg  _T_344; // @[Reg.scala 15:16]
  reg  _T_345; // @[Reg.scala 15:16]
  reg  _T_346; // @[Reg.scala 15:16]
  reg  _T_347; // @[Reg.scala 15:16]
  reg  _T_348; // @[Reg.scala 15:16]
  reg  _T_349; // @[Reg.scala 15:16]
  reg  _T_350; // @[Reg.scala 15:16]
  reg  _T_351; // @[Reg.scala 15:16]
  reg  _T_352; // @[Reg.scala 15:16]
  reg  _T_353; // @[Reg.scala 15:16]
  reg  _T_354; // @[Reg.scala 15:16]
  reg  _T_355; // @[Reg.scala 15:16]
  reg  _T_356; // @[Reg.scala 15:16]
  reg  _T_357; // @[Reg.scala 15:16]
  reg  _T_358; // @[Reg.scala 15:16]
  reg  _T_359; // @[Reg.scala 15:16]
  reg  _T_360; // @[Reg.scala 15:16]
  reg  _T_361; // @[Reg.scala 15:16]
  reg  _T_362; // @[Reg.scala 15:16]
  reg  _T_363; // @[Reg.scala 15:16]
  reg  _T_364; // @[Reg.scala 15:16]
  reg  _T_365; // @[Reg.scala 15:16]
  reg  _T_366; // @[Reg.scala 15:16]
  reg  _T_367; // @[Reg.scala 15:16]
  reg  _T_368; // @[Reg.scala 15:16]
  reg  _T_369; // @[Reg.scala 15:16]
  reg  _T_370; // @[Reg.scala 15:16]
  reg  _T_371; // @[Reg.scala 15:16]
  reg  _T_372; // @[Reg.scala 15:16]
  reg  _T_373; // @[Reg.scala 15:16]
  reg  _T_374; // @[Reg.scala 15:16]
  reg  _T_375; // @[Reg.scala 15:16]
  reg  _T_376; // @[Reg.scala 15:16]
  reg  _T_377; // @[Reg.scala 15:16]
  reg  _T_378; // @[Reg.scala 15:16]
  reg  _T_379; // @[Reg.scala 15:16]
  reg  _T_380; // @[Reg.scala 15:16]
  reg  _T_381; // @[Reg.scala 15:16]
  reg  _T_382; // @[Reg.scala 15:16]
  reg  _T_383; // @[Reg.scala 15:16]
  reg  _T_384; // @[Reg.scala 15:16]
  reg  _T_385; // @[Reg.scala 15:16]
  reg  _T_386; // @[Reg.scala 15:16]
  reg  _T_387; // @[Reg.scala 15:16]
  reg  _T_388; // @[Reg.scala 15:16]
  reg  _T_389; // @[Reg.scala 15:16]
  reg  _T_390; // @[Reg.scala 15:16]
  reg  _T_391; // @[Reg.scala 15:16]
  reg  _T_392; // @[Reg.scala 15:16]
  reg  _T_393; // @[Reg.scala 15:16]
  reg  _T_394; // @[Reg.scala 15:16]
  reg  _T_395; // @[Reg.scala 15:16]
  reg  _T_396; // @[Reg.scala 15:16]
  reg  _T_397; // @[Reg.scala 15:16]
  reg  _T_398; // @[Reg.scala 15:16]
  reg  _T_399; // @[Reg.scala 15:16]
  reg  _T_400; // @[Reg.scala 15:16]
  reg  _T_401; // @[Reg.scala 15:16]
  reg  _T_402; // @[Reg.scala 15:16]
  reg  _T_403; // @[Reg.scala 15:16]
  reg  _T_404; // @[Reg.scala 15:16]
  reg  _T_405; // @[Reg.scala 15:16]
  reg  _T_406; // @[Reg.scala 15:16]
  reg  _T_407; // @[Reg.scala 15:16]
  reg  _T_408; // @[Reg.scala 15:16]
  reg  _T_409; // @[Reg.scala 15:16]
  reg  _T_410; // @[Reg.scala 15:16]
  reg  _T_411; // @[Reg.scala 15:16]
  reg  _T_412; // @[Reg.scala 15:16]
  reg  _T_413; // @[Reg.scala 15:16]
  reg  _T_414; // @[Reg.scala 15:16]
  reg  _T_415; // @[Reg.scala 15:16]
  reg  _T_416; // @[Reg.scala 15:16]
  reg  _T_417; // @[Reg.scala 15:16]
  reg  _T_418; // @[Reg.scala 15:16]
  reg  _T_419; // @[Reg.scala 15:16]
  reg  _T_420; // @[Reg.scala 15:16]
  reg  _T_421; // @[Reg.scala 15:16]
  reg  _T_422; // @[Reg.scala 15:16]
  reg  _T_423; // @[Reg.scala 15:16]
  reg  _T_424; // @[Reg.scala 15:16]
  reg  _T_425; // @[Reg.scala 15:16]
  reg  _T_426; // @[Reg.scala 15:16]
  reg  _T_427; // @[Reg.scala 15:16]
  reg  _T_428; // @[Reg.scala 15:16]
  reg  _T_429; // @[Reg.scala 15:16]
  reg  _T_430; // @[Reg.scala 15:16]
  reg  _T_431; // @[Reg.scala 15:16]
  reg  _T_432; // @[Reg.scala 15:16]
  reg  _T_433; // @[Reg.scala 15:16]
  reg  _T_434; // @[Reg.scala 15:16]
  reg  _T_435; // @[Reg.scala 15:16]
  reg  _T_436; // @[Reg.scala 15:16]
  reg  _T_437; // @[Reg.scala 15:16]
  reg  _T_438; // @[Reg.scala 15:16]
  reg  _T_439; // @[Reg.scala 15:16]
  reg  _T_440; // @[Reg.scala 15:16]
  reg  _T_441; // @[Reg.scala 15:16]
  reg  _T_442; // @[Reg.scala 15:16]
  reg  _T_443; // @[Reg.scala 15:16]
  reg  _T_444; // @[Reg.scala 15:16]
  reg  _T_445; // @[Reg.scala 15:16]
  reg  _T_446; // @[Reg.scala 15:16]
  reg  _T_447; // @[Reg.scala 15:16]
  reg  _T_448; // @[Reg.scala 15:16]
  reg  _T_449; // @[Reg.scala 15:16]
  reg  _T_450; // @[Reg.scala 15:16]
  reg  _T_451; // @[Reg.scala 15:16]
  reg  _T_452; // @[Reg.scala 15:16]
  reg  _T_453; // @[Reg.scala 15:16]
  reg  _T_454; // @[Reg.scala 15:16]
  reg  _T_455; // @[Reg.scala 15:16]
  reg  _T_456; // @[Reg.scala 15:16]
  reg  _T_457; // @[Reg.scala 15:16]
  reg  _T_458; // @[Reg.scala 15:16]
  reg  _T_459; // @[Reg.scala 15:16]
  reg  _T_460; // @[Reg.scala 15:16]
  reg  _T_461; // @[Reg.scala 15:16]
  reg  _T_462; // @[Reg.scala 15:16]
  reg  _T_463; // @[Reg.scala 15:16]
  reg  _T_464; // @[Reg.scala 15:16]
  reg  _T_465; // @[Reg.scala 15:16]
  reg  _T_466; // @[Reg.scala 15:16]
  reg  _T_467; // @[Reg.scala 15:16]
  reg  _T_468; // @[Reg.scala 15:16]
  reg  _T_469; // @[Reg.scala 15:16]
  reg  _T_470; // @[Reg.scala 15:16]
  reg  _T_471; // @[Reg.scala 15:16]
  reg  _T_472; // @[Reg.scala 15:16]
  reg  _T_473; // @[Reg.scala 15:16]
  reg  _T_474; // @[Reg.scala 15:16]
  reg  _T_475; // @[Reg.scala 15:16]
  reg  _T_476; // @[Reg.scala 15:16]
  reg  _T_477; // @[Reg.scala 15:16]
  reg  _T_478; // @[Reg.scala 15:16]
  reg  _T_479; // @[Reg.scala 15:16]
  reg  _T_480; // @[Reg.scala 15:16]
  reg  _T_481; // @[Reg.scala 15:16]
  reg  _T_482; // @[Reg.scala 15:16]
  reg  _T_483; // @[Reg.scala 15:16]
  reg  _T_484; // @[Reg.scala 15:16]
  reg  _T_485; // @[Reg.scala 15:16]
  reg  _T_486; // @[Reg.scala 15:16]
  reg  _T_487; // @[Reg.scala 15:16]
  reg  _T_488; // @[Reg.scala 15:16]
  reg  _T_489; // @[Reg.scala 15:16]
  reg  _T_490; // @[Reg.scala 15:16]
  reg  _T_491; // @[Reg.scala 15:16]
  reg  _T_492; // @[Reg.scala 15:16]
  reg  _T_493; // @[Reg.scala 15:16]
  reg  _T_494; // @[Reg.scala 15:16]
  reg  _T_495; // @[Reg.scala 15:16]
  reg  _T_496; // @[Reg.scala 15:16]
  reg  _T_497; // @[Reg.scala 15:16]
  reg  _T_498; // @[Reg.scala 15:16]
  reg  _T_499; // @[Reg.scala 15:16]
  reg  _T_500; // @[Reg.scala 15:16]
  reg  _T_501; // @[Reg.scala 15:16]
  reg  _T_502; // @[Reg.scala 15:16]
  reg  _T_503; // @[Reg.scala 15:16]
  reg  _T_504; // @[Reg.scala 15:16]
  reg  _T_505; // @[Reg.scala 15:16]
  reg  _T_506; // @[Reg.scala 15:16]
  reg  _T_507; // @[Reg.scala 15:16]
  reg  _T_508; // @[Reg.scala 15:16]
  reg  _T_509; // @[Reg.scala 15:16]
  reg  _T_510; // @[Reg.scala 15:16]
  reg  _T_511; // @[Reg.scala 15:16]
  reg  _T_512; // @[Reg.scala 15:16]
  reg  _T_513; // @[Reg.scala 15:16]
  reg  _T_514; // @[Reg.scala 15:16]
  reg  _T_515; // @[Reg.scala 15:16]
  reg  _T_516; // @[Reg.scala 15:16]
  reg  _T_517; // @[Reg.scala 15:16]
  reg  _T_518; // @[Reg.scala 15:16]
  reg  _T_519; // @[Reg.scala 15:16]
  reg  _T_520; // @[Reg.scala 15:16]
  reg  _T_521; // @[Reg.scala 15:16]
  reg  _T_522; // @[Reg.scala 15:16]
  reg  _T_523; // @[Reg.scala 15:16]
  reg  _T_524; // @[Reg.scala 15:16]
  reg  _T_525; // @[Reg.scala 15:16]
  reg  _T_526; // @[Reg.scala 15:16]
  reg  _T_527; // @[Reg.scala 15:16]
  reg  _T_528; // @[Reg.scala 15:16]
  reg  _T_529; // @[Reg.scala 15:16]
  reg  _T_530; // @[Reg.scala 15:16]
  reg  _T_531; // @[Reg.scala 15:16]
  reg  _T_532; // @[Reg.scala 15:16]
  reg  _T_533; // @[Reg.scala 15:16]
  reg  _T_534; // @[Reg.scala 15:16]
  reg  _T_535; // @[Reg.scala 15:16]
  reg  _T_536; // @[Reg.scala 15:16]
  reg  _T_537; // @[Reg.scala 15:16]
  reg  _T_538; // @[Reg.scala 15:16]
  reg  _T_539; // @[Reg.scala 15:16]
  reg  _T_540; // @[Reg.scala 15:16]
  reg  _T_541; // @[Reg.scala 15:16]
  reg  _T_542; // @[Reg.scala 15:16]
  reg  _T_543; // @[Reg.scala 15:16]
  reg  _T_544; // @[Reg.scala 15:16]
  reg  _T_545; // @[Reg.scala 15:16]
  reg  _T_546; // @[Reg.scala 15:16]
  reg  _T_547; // @[Reg.scala 15:16]
  reg  _T_548; // @[Reg.scala 15:16]
  reg  _T_549; // @[Reg.scala 15:16]
  reg  _T_550; // @[Reg.scala 15:16]
  reg  _T_551; // @[Reg.scala 15:16]
  reg  _T_552; // @[Reg.scala 15:16]
  reg  _T_553; // @[Reg.scala 15:16]
  reg  _T_554; // @[Reg.scala 15:16]
  reg  _T_555; // @[Reg.scala 15:16]
  reg  _T_556; // @[Reg.scala 15:16]
  reg  _T_557; // @[Reg.scala 15:16]
  reg  _T_558; // @[Reg.scala 15:16]
  reg  _T_559; // @[Reg.scala 15:16]
  reg  _T_560; // @[Reg.scala 15:16]
  reg  _T_561; // @[Reg.scala 15:16]
  reg  _T_562; // @[Reg.scala 15:16]
  reg  _T_563; // @[Reg.scala 15:16]
  reg  _T_564; // @[Reg.scala 15:16]
  reg  _T_565; // @[Reg.scala 15:16]
  reg  _T_566; // @[Reg.scala 15:16]
  reg  _T_567; // @[Reg.scala 15:16]
  reg  _T_568; // @[Reg.scala 15:16]
  reg  _T_569; // @[Reg.scala 15:16]
  reg  _T_570; // @[Reg.scala 15:16]
  reg  _T_571; // @[Reg.scala 15:16]
  reg  _T_572; // @[Reg.scala 15:16]
  reg  _T_573; // @[Reg.scala 15:16]
  reg  _T_574; // @[Reg.scala 15:16]
  reg  _T_575; // @[Reg.scala 15:16]
  reg  _T_576; // @[Reg.scala 15:16]
  reg  _T_577; // @[Reg.scala 15:16]
  reg  _T_578; // @[Reg.scala 15:16]
  reg  _T_579; // @[Reg.scala 15:16]
  reg  _T_580; // @[Reg.scala 15:16]
  reg  _T_581; // @[Reg.scala 15:16]
  reg  _T_582; // @[Reg.scala 15:16]
  reg  _T_583; // @[Reg.scala 15:16]
  reg  _T_584; // @[Reg.scala 15:16]
  reg  _T_585; // @[Reg.scala 15:16]
  reg  _T_586; // @[Reg.scala 15:16]
  reg  _T_587; // @[Reg.scala 15:16]
  reg  _T_588; // @[Reg.scala 15:16]
  reg  _T_589; // @[Reg.scala 15:16]
  reg  _T_590; // @[Reg.scala 15:16]
  reg  _T_591; // @[Reg.scala 15:16]
  reg  _T_592; // @[Reg.scala 15:16]
  reg  _T_593; // @[Reg.scala 15:16]
  reg  _T_594; // @[Reg.scala 15:16]
  reg  _T_595; // @[Reg.scala 15:16]
  reg  _T_596; // @[Reg.scala 15:16]
  reg  _T_597; // @[Reg.scala 15:16]
  reg  _T_598; // @[Reg.scala 15:16]
  reg  _T_599; // @[Reg.scala 15:16]
  reg  _T_600; // @[Reg.scala 15:16]
  reg  _T_601; // @[Reg.scala 15:16]
  reg  _T_602; // @[Reg.scala 15:16]
  reg  _T_603; // @[Reg.scala 15:16]
  reg  _T_604; // @[Reg.scala 15:16]
  reg  _T_605; // @[Reg.scala 15:16]
  reg  _T_606; // @[Reg.scala 15:16]
  reg  _T_607; // @[Reg.scala 15:16]
  reg  _T_608; // @[Reg.scala 15:16]
  reg  _T_609; // @[Reg.scala 15:16]
  reg  _T_610; // @[Reg.scala 15:16]
  reg  _T_611; // @[Reg.scala 15:16]
  reg  _T_612; // @[Reg.scala 15:16]
  reg  _T_613; // @[Reg.scala 15:16]
  reg  _T_614; // @[Reg.scala 15:16]
  reg  _T_615; // @[Reg.scala 15:16]
  reg  _T_616; // @[Reg.scala 15:16]
  reg  _T_617; // @[Reg.scala 15:16]
  reg  _T_618; // @[Reg.scala 15:16]
  reg  _T_619; // @[Reg.scala 15:16]
  reg  _T_620; // @[Reg.scala 15:16]
  reg  _T_621; // @[Reg.scala 15:16]
  reg  _T_622; // @[Reg.scala 15:16]
  reg  _T_623; // @[Reg.scala 15:16]
  reg  _T_624; // @[Reg.scala 15:16]
  reg  _T_625; // @[Reg.scala 15:16]
  reg  _T_626; // @[Reg.scala 15:16]
  reg  _T_627; // @[Reg.scala 15:16]
  reg  _T_628; // @[Reg.scala 15:16]
  reg  _T_629; // @[Reg.scala 15:16]
  reg  _T_630; // @[Reg.scala 15:16]
  reg  _T_631; // @[Reg.scala 15:16]
  reg  _T_632; // @[Reg.scala 15:16]
  reg  _T_633; // @[Reg.scala 15:16]
  reg  _T_634; // @[Reg.scala 15:16]
  reg  _T_635; // @[Reg.scala 15:16]
  reg  _T_636; // @[Reg.scala 15:16]
  reg  _T_637; // @[Reg.scala 15:16]
  reg  _T_638; // @[Reg.scala 15:16]
  reg  _T_639; // @[Reg.scala 15:16]
  reg  _T_640; // @[Reg.scala 15:16]
  reg  _T_641; // @[Reg.scala 15:16]
  reg  _T_642; // @[Reg.scala 15:16]
  reg  _T_643; // @[Reg.scala 15:16]
  reg  _T_644; // @[Reg.scala 15:16]
  reg  _T_645; // @[Reg.scala 15:16]
  reg  _T_646; // @[Reg.scala 15:16]
  reg  _T_647; // @[Reg.scala 15:16]
  reg  _T_648; // @[Reg.scala 15:16]
  reg  _T_649; // @[Reg.scala 15:16]
  reg  _T_650; // @[Reg.scala 15:16]
  reg  _T_651; // @[Reg.scala 15:16]
  reg  _T_652; // @[Reg.scala 15:16]
  reg  _T_653; // @[Reg.scala 15:16]
  reg  _T_654; // @[Reg.scala 15:16]
  reg  _T_655; // @[Reg.scala 15:16]
  reg  _T_656; // @[Reg.scala 15:16]
  reg  _T_657; // @[Reg.scala 15:16]
  reg  _T_658; // @[Reg.scala 15:16]
  reg  _T_659; // @[Reg.scala 15:16]
  reg  _T_660; // @[Reg.scala 15:16]
  reg  _T_661; // @[Reg.scala 15:16]
  reg  _T_662; // @[Reg.scala 15:16]
  reg  _T_663; // @[Reg.scala 15:16]
  reg  _T_664; // @[Reg.scala 15:16]
  reg  _T_665; // @[Reg.scala 15:16]
  reg  _T_666; // @[Reg.scala 15:16]
  reg  _T_667; // @[Reg.scala 15:16]
  reg  _T_668; // @[Reg.scala 15:16]
  reg  _T_669; // @[Reg.scala 15:16]
  reg  _T_670; // @[Reg.scala 15:16]
  reg  _T_671; // @[Reg.scala 15:16]
  reg  _T_672; // @[Reg.scala 15:16]
  reg  _T_673; // @[Reg.scala 15:16]
  reg  _T_674; // @[Reg.scala 15:16]
  reg  _T_675; // @[Reg.scala 15:16]
  reg  _T_676; // @[Reg.scala 15:16]
  reg  _T_677; // @[Reg.scala 15:16]
  reg  _T_678; // @[Reg.scala 15:16]
  reg  _T_679; // @[Reg.scala 15:16]
  reg  _T_680; // @[Reg.scala 15:16]
  reg  _T_681; // @[Reg.scala 15:16]
  reg  _T_682; // @[Reg.scala 15:16]
  reg  _T_683; // @[Reg.scala 15:16]
  reg  _T_684; // @[Reg.scala 15:16]
  reg  _T_685; // @[Reg.scala 15:16]
  reg  _T_686; // @[Reg.scala 15:16]
  reg  _T_687; // @[Reg.scala 15:16]
  reg  _T_688; // @[Reg.scala 15:16]
  reg  _T_689; // @[Reg.scala 15:16]
  reg  _T_690; // @[Reg.scala 15:16]
  reg  _T_691; // @[Reg.scala 15:16]
  reg  _T_692; // @[Reg.scala 15:16]
  reg  _T_693; // @[Reg.scala 15:16]
  reg  _T_694; // @[Reg.scala 15:16]
  reg  _T_695; // @[Reg.scala 15:16]
  reg  _T_696; // @[Reg.scala 15:16]
  reg  _T_697; // @[Reg.scala 15:16]
  reg  _T_698; // @[Reg.scala 15:16]
  reg  _T_699; // @[Reg.scala 15:16]
  reg  _T_700; // @[Reg.scala 15:16]
  reg  _T_701; // @[Reg.scala 15:16]
  reg  _T_702; // @[Reg.scala 15:16]
  reg  _T_703; // @[Reg.scala 15:16]
  reg  _T_704; // @[Reg.scala 15:16]
  reg  _T_705; // @[Reg.scala 15:16]
  reg  _T_706; // @[Reg.scala 15:16]
  reg  _T_707; // @[Reg.scala 15:16]
  reg  _T_708; // @[Reg.scala 15:16]
  reg  _T_709; // @[Reg.scala 15:16]
  reg  _T_710; // @[Reg.scala 15:16]
  reg  _T_711; // @[Reg.scala 15:16]
  reg  _T_712; // @[Reg.scala 15:16]
  reg  _T_713; // @[Reg.scala 15:16]
  reg  _T_714; // @[Reg.scala 15:16]
  reg  _T_715; // @[Reg.scala 15:16]
  reg  _T_716; // @[Reg.scala 15:16]
  reg  _T_717; // @[Reg.scala 15:16]
  reg  _T_718; // @[Reg.scala 15:16]
  reg  _T_719; // @[Reg.scala 15:16]
  reg  _T_720; // @[Reg.scala 15:16]
  reg  _T_721; // @[Reg.scala 15:16]
  reg  _T_722; // @[Reg.scala 15:16]
  reg  _T_723; // @[Reg.scala 15:16]
  reg  _T_724; // @[Reg.scala 15:16]
  reg  _T_725; // @[Reg.scala 15:16]
  reg  _T_726; // @[Reg.scala 15:16]
  reg  _T_727; // @[Reg.scala 15:16]
  reg  _T_728; // @[Reg.scala 15:16]
  reg  _T_729; // @[Reg.scala 15:16]
  reg  _T_730; // @[Reg.scala 15:16]
  reg  _T_731; // @[Reg.scala 15:16]
  reg  _T_732; // @[Reg.scala 15:16]
  reg  _T_733; // @[Reg.scala 15:16]
  reg  _T_734; // @[Reg.scala 15:16]
  reg  _T_735; // @[Reg.scala 15:16]
  reg  _T_736; // @[Reg.scala 15:16]
  reg  _T_737; // @[Reg.scala 15:16]
  reg  _T_738; // @[Reg.scala 15:16]
  reg  _T_739; // @[Reg.scala 15:16]
  reg  _T_740; // @[Reg.scala 15:16]
  reg  _T_741; // @[Reg.scala 15:16]
  reg  _T_742; // @[Reg.scala 15:16]
  reg  _T_743; // @[Reg.scala 15:16]
  reg  _T_744; // @[Reg.scala 15:16]
  reg  _T_745; // @[Reg.scala 15:16]
  reg  _T_746; // @[Reg.scala 15:16]
  reg  _T_747; // @[Reg.scala 15:16]
  reg  _T_748; // @[Reg.scala 15:16]
  reg  _T_749; // @[Reg.scala 15:16]
  reg  _T_750; // @[Reg.scala 15:16]
  reg  _T_751; // @[Reg.scala 15:16]
  reg  _T_752; // @[Reg.scala 15:16]
  reg  _T_753; // @[Reg.scala 15:16]
  reg  _T_754; // @[Reg.scala 15:16]
  reg  _T_755; // @[Reg.scala 15:16]
  reg  _T_756; // @[Reg.scala 15:16]
  reg  _T_757; // @[Reg.scala 15:16]
  reg  _T_758; // @[Reg.scala 15:16]
  reg  _T_759; // @[Reg.scala 15:16]
  reg  _T_760; // @[Reg.scala 15:16]
  reg  _T_761; // @[Reg.scala 15:16]
  reg  _T_762; // @[Reg.scala 15:16]
  reg  _T_763; // @[Reg.scala 15:16]
  reg  _T_764; // @[Reg.scala 15:16]
  reg  _T_765; // @[Reg.scala 15:16]
  reg  _T_766; // @[Reg.scala 15:16]
  reg  _T_767; // @[Reg.scala 15:16]
  reg  _T_768; // @[Reg.scala 15:16]
  reg  _T_769; // @[Reg.scala 15:16]
  reg  _T_770; // @[Reg.scala 15:16]
  reg  _T_771; // @[Reg.scala 15:16]
  reg  _T_772; // @[Reg.scala 15:16]
  reg  _T_773; // @[Reg.scala 15:16]
  reg  _T_774; // @[Reg.scala 15:16]
  reg  _T_775; // @[Reg.scala 15:16]
  reg  _T_776; // @[Reg.scala 15:16]
  reg  _T_777; // @[Reg.scala 15:16]
  reg  _T_778; // @[Reg.scala 15:16]
  reg  _T_779; // @[Reg.scala 15:16]
  reg  _T_780; // @[Reg.scala 15:16]
  reg  _T_781; // @[Reg.scala 15:16]
  reg  _T_782; // @[Reg.scala 15:16]
  reg  _T_783; // @[Reg.scala 15:16]
  reg  _T_784; // @[Reg.scala 15:16]
  reg  _T_785; // @[Reg.scala 15:16]
  reg  _T_786; // @[Reg.scala 15:16]
  reg  _T_787; // @[Reg.scala 15:16]
  reg  _T_788; // @[Reg.scala 15:16]
  reg  _T_789; // @[Reg.scala 15:16]
  reg  _T_790; // @[Reg.scala 15:16]
  reg  _T_791; // @[Reg.scala 15:16]
  reg  _T_792; // @[Reg.scala 15:16]
  reg  _T_793; // @[Reg.scala 15:16]
  reg  _T_794; // @[Reg.scala 15:16]
  reg  _T_795; // @[Reg.scala 15:16]
  reg  _T_796; // @[Reg.scala 15:16]
  reg  _T_797; // @[Reg.scala 15:16]
  reg  _T_798; // @[Reg.scala 15:16]
  reg  _T_799; // @[Reg.scala 15:16]
  reg  _T_800; // @[Reg.scala 15:16]
  reg  _T_801; // @[Reg.scala 15:16]
  reg  _T_802; // @[Reg.scala 15:16]
  reg  _T_803; // @[Reg.scala 15:16]
  reg  _T_804; // @[Reg.scala 15:16]
  reg  _T_805; // @[Reg.scala 15:16]
  reg  _T_806; // @[Reg.scala 15:16]
  reg  _T_807; // @[Reg.scala 15:16]
  reg  _T_808; // @[Reg.scala 15:16]
  reg  _T_809; // @[Reg.scala 15:16]
  reg  _T_810; // @[Reg.scala 15:16]
  reg  _T_811; // @[Reg.scala 15:16]
  reg  _T_812; // @[Reg.scala 15:16]
  reg  _T_813; // @[Reg.scala 15:16]
  reg  _T_814; // @[Reg.scala 15:16]
  reg  _T_815; // @[Reg.scala 15:16]
  reg  _T_816; // @[Reg.scala 15:16]
  reg  _T_817; // @[Reg.scala 15:16]
  reg  _T_818; // @[Reg.scala 15:16]
  reg  _T_819; // @[Reg.scala 15:16]
  reg  _T_820; // @[Reg.scala 15:16]
  reg  _T_821; // @[Reg.scala 15:16]
  reg  _T_822; // @[Reg.scala 15:16]
  reg  _T_823; // @[Reg.scala 15:16]
  reg  _T_824; // @[Reg.scala 15:16]
  reg  _T_825; // @[Reg.scala 15:16]
  reg  _T_826; // @[Reg.scala 15:16]
  reg  _T_827; // @[Reg.scala 15:16]
  reg  _T_828; // @[Reg.scala 15:16]
  reg  _T_829; // @[Reg.scala 15:16]
  reg  _T_830; // @[Reg.scala 15:16]
  reg  _T_831; // @[Reg.scala 15:16]
  reg  _T_832; // @[Reg.scala 15:16]
  reg  _T_833; // @[Reg.scala 15:16]
  reg  _T_834; // @[Reg.scala 15:16]
  reg  _T_835; // @[Reg.scala 15:16]
  reg  _T_836; // @[Reg.scala 15:16]
  reg  _T_837; // @[Reg.scala 15:16]
  reg  _T_838; // @[Reg.scala 15:16]
  reg  _T_839; // @[Reg.scala 15:16]
  wire [8:0] _T_842 = out_counter + 9'h1; // @[Reorder.scala 41:32]
  wire  _T_843 = out_counter < 9'h100; // @[Reorder.scala 44:20]
  assign rambank0_re__T_845_addr = out_counter[7:0];
  assign rambank0_re__T_845_data = rambank0_re[rambank0_re__T_845_addr]; // @[Reorder.scala 20:21]
  assign rambank0_re__T_69_data = io_in1_re;
  assign rambank0_re__T_69_addr = index1[7:0];
  assign rambank0_re__T_69_mask = 1'h1;
  assign rambank0_re__T_69_en = io_in_valid & _T_64;
  assign rambank0_im__T_845_addr = out_counter[7:0];
  assign rambank0_im__T_845_data = rambank0_im[rambank0_im__T_845_addr]; // @[Reorder.scala 20:21]
  assign rambank0_im__T_69_data = io_in1_im;
  assign rambank0_im__T_69_addr = index1[7:0];
  assign rambank0_im__T_69_mask = 1'h1;
  assign rambank0_im__T_69_en = io_in_valid & _T_64;
  assign rambank1_re__T_847_addr = out_counter[7:0];
  assign rambank1_re__T_847_data = rambank1_re[rambank1_re__T_847_addr]; // @[Reorder.scala 21:21]
  assign rambank1_re__T_71_data = io_in2_re;
  assign rambank1_re__T_71_addr = index2[7:0];
  assign rambank1_re__T_71_mask = 1'h1;
  assign rambank1_re__T_71_en = io_in_valid & _T_64;
  assign rambank1_im__T_847_addr = out_counter[7:0];
  assign rambank1_im__T_847_data = rambank1_im[rambank1_im__T_847_addr]; // @[Reorder.scala 21:21]
  assign rambank1_im__T_71_data = io_in2_im;
  assign rambank1_im__T_71_addr = index2[7:0];
  assign rambank1_im__T_71_mask = 1'h1;
  assign rambank1_im__T_71_en = io_in_valid & _T_64;
  assign io_out_re = _T_843 ? $signed(rambank0_re__T_845_data) : $signed(rambank1_re__T_847_data); // @[Reorder.scala 45:12 Reorder.scala 47:12]
  assign io_out_im = _T_843 ? $signed(rambank0_im__T_845_data) : $signed(rambank1_im__T_847_data); // @[Reorder.scala 45:12 Reorder.scala 47:12]
  assign io_out_valid = _T_327 | _T_839; // @[Reorder.scala 39:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank0_re[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank0_im[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank1_re[initvar] = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    rambank1_im[initvar] = _RAND_3[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_counter = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  out_counter = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  _T_72 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_73 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_74 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_75 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_76 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_77 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_78 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_79 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_80 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_81 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_82 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_83 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_84 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_85 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_86 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_87 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_88 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_89 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_90 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_91 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  _T_92 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_93 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  _T_94 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_95 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  _T_96 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_97 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_98 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_99 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_100 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_101 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_102 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_103 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_104 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_105 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_106 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_107 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_108 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_109 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_110 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_111 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_112 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_113 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  _T_114 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_115 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_116 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_117 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  _T_118 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  _T_119 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  _T_120 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  _T_121 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_122 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  _T_123 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  _T_124 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  _T_125 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  _T_126 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  _T_127 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_128 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_129 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_130 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_131 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _T_132 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  _T_133 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _T_134 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _T_135 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _T_136 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _T_137 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _T_138 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _T_139 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _T_140 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  _T_141 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _T_142 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  _T_143 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  _T_144 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  _T_145 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  _T_146 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  _T_147 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  _T_148 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  _T_149 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  _T_150 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  _T_151 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  _T_152 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  _T_153 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  _T_154 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  _T_155 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  _T_156 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  _T_157 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  _T_158 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _T_159 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_160 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _T_161 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _T_162 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _T_163 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _T_164 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _T_165 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _T_166 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  _T_167 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  _T_168 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  _T_169 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  _T_170 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _T_171 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  _T_172 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  _T_173 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _T_174 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  _T_175 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  _T_176 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  _T_177 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  _T_178 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  _T_179 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  _T_180 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  _T_181 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  _T_182 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  _T_183 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  _T_184 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  _T_185 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  _T_186 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  _T_187 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  _T_188 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  _T_189 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  _T_190 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  _T_191 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  _T_192 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  _T_193 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  _T_194 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  _T_195 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  _T_196 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  _T_197 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  _T_198 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  _T_199 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  _T_200 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  _T_201 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  _T_202 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  _T_203 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  _T_204 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  _T_205 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  _T_206 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  _T_207 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  _T_208 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  _T_209 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  _T_210 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  _T_211 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  _T_212 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  _T_213 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  _T_214 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  _T_215 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  _T_216 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  _T_217 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  _T_218 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  _T_219 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  _T_220 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  _T_221 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  _T_222 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  _T_223 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  _T_224 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  _T_225 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  _T_226 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  _T_227 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  _T_228 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  _T_229 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  _T_230 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  _T_231 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  _T_232 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  _T_233 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  _T_234 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  _T_235 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  _T_236 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  _T_237 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  _T_238 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  _T_239 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  _T_240 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  _T_241 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  _T_242 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  _T_243 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  _T_244 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  _T_245 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  _T_246 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  _T_247 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  _T_248 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  _T_249 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  _T_250 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  _T_251 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  _T_252 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  _T_253 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  _T_254 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  _T_255 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  _T_256 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  _T_257 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  _T_258 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  _T_259 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  _T_260 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  _T_261 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  _T_262 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  _T_263 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  _T_264 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  _T_265 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  _T_266 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  _T_267 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  _T_268 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  _T_269 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  _T_270 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  _T_271 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  _T_272 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  _T_273 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  _T_274 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  _T_275 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  _T_276 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  _T_277 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  _T_278 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  _T_279 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  _T_280 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  _T_281 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  _T_282 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  _T_283 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  _T_284 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  _T_285 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  _T_286 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  _T_287 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  _T_288 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  _T_289 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  _T_290 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  _T_291 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  _T_292 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  _T_293 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  _T_294 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  _T_295 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  _T_296 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  _T_297 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  _T_298 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  _T_299 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  _T_300 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  _T_301 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  _T_302 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  _T_303 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  _T_304 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  _T_305 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  _T_306 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  _T_307 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  _T_308 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  _T_309 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  _T_310 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  _T_311 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  _T_312 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  _T_313 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  _T_314 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  _T_315 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  _T_316 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  _T_317 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  _T_318 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  _T_319 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  _T_320 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  _T_321 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  _T_322 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  _T_323 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  _T_324 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  _T_325 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  _T_326 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  _T_327 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  _T_328 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  _T_329 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  _T_330 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  _T_331 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  _T_332 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  _T_333 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  _T_334 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  _T_335 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  _T_336 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  _T_337 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  _T_338 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  _T_339 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  _T_340 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  _T_341 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  _T_342 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  _T_343 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  _T_344 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  _T_345 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  _T_346 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  _T_347 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  _T_348 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  _T_349 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  _T_350 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  _T_351 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  _T_352 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  _T_353 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  _T_354 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  _T_355 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  _T_356 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  _T_357 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  _T_358 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  _T_359 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  _T_360 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  _T_361 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  _T_362 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  _T_363 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  _T_364 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  _T_365 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  _T_366 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  _T_367 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  _T_368 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  _T_369 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  _T_370 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  _T_371 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  _T_372 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  _T_373 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  _T_374 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  _T_375 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  _T_376 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  _T_377 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  _T_378 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  _T_379 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  _T_380 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  _T_381 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  _T_382 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  _T_383 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  _T_384 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  _T_385 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  _T_386 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  _T_387 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  _T_388 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  _T_389 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  _T_390 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  _T_391 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  _T_392 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  _T_393 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  _T_394 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  _T_395 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  _T_396 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  _T_397 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  _T_398 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  _T_399 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  _T_400 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  _T_401 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  _T_402 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  _T_403 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  _T_404 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  _T_405 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  _T_406 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  _T_407 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  _T_408 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  _T_409 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  _T_410 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  _T_411 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  _T_412 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  _T_413 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  _T_414 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  _T_415 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  _T_416 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  _T_417 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  _T_418 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  _T_419 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  _T_420 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  _T_421 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  _T_422 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  _T_423 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  _T_424 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  _T_425 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  _T_426 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  _T_427 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  _T_428 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  _T_429 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  _T_430 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  _T_431 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  _T_432 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  _T_433 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  _T_434 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  _T_435 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  _T_436 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  _T_437 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  _T_438 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  _T_439 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  _T_440 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  _T_441 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  _T_442 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  _T_443 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  _T_444 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  _T_445 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  _T_446 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  _T_447 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  _T_448 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  _T_449 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  _T_450 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  _T_451 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  _T_452 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  _T_453 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  _T_454 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  _T_455 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  _T_456 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  _T_457 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  _T_458 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  _T_459 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  _T_460 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  _T_461 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  _T_462 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  _T_463 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  _T_464 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  _T_465 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  _T_466 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  _T_467 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  _T_468 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  _T_469 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  _T_470 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  _T_471 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  _T_472 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  _T_473 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  _T_474 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  _T_475 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  _T_476 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  _T_477 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  _T_478 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  _T_479 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  _T_480 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  _T_481 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  _T_482 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  _T_483 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  _T_484 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  _T_485 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  _T_486 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  _T_487 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  _T_488 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  _T_489 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  _T_490 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  _T_491 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  _T_492 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  _T_493 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  _T_494 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  _T_495 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  _T_496 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  _T_497 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  _T_498 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  _T_499 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  _T_500 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  _T_501 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  _T_502 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  _T_503 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  _T_504 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  _T_505 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  _T_506 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  _T_507 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  _T_508 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  _T_509 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  _T_510 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  _T_511 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  _T_512 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  _T_513 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  _T_514 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  _T_515 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  _T_516 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  _T_517 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  _T_518 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  _T_519 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  _T_520 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  _T_521 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  _T_522 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  _T_523 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  _T_524 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  _T_525 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  _T_526 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  _T_527 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  _T_528 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_529 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_530 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_531 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_532 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_533 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_534 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_535 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_536 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_537 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_538 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  _T_539 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  _T_540 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  _T_541 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  _T_542 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  _T_543 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  _T_544 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  _T_545 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  _T_546 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  _T_547 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  _T_548 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  _T_549 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  _T_550 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  _T_551 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  _T_552 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  _T_553 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  _T_554 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  _T_555 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  _T_556 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  _T_557 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  _T_558 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  _T_559 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  _T_560 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  _T_561 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  _T_562 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  _T_563 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  _T_564 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  _T_565 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  _T_566 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  _T_567 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  _T_568 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  _T_569 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  _T_570 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  _T_571 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  _T_572 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  _T_573 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  _T_574 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  _T_575 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  _T_576 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  _T_577 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  _T_578 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  _T_579 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  _T_580 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  _T_581 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  _T_582 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  _T_583 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  _T_584 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  _T_585 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  _T_586 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  _T_587 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  _T_588 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  _T_589 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  _T_590 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  _T_591 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  _T_592 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  _T_593 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  _T_594 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  _T_595 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  _T_596 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  _T_597 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  _T_598 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  _T_599 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  _T_600 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  _T_601 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  _T_602 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  _T_603 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  _T_604 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  _T_605 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  _T_606 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  _T_607 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  _T_608 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  _T_609 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  _T_610 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  _T_611 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  _T_612 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  _T_613 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  _T_614 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  _T_615 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  _T_616 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  _T_617 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  _T_618 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  _T_619 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  _T_620 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  _T_621 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  _T_622 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  _T_623 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  _T_624 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  _T_625 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  _T_626 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  _T_627 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  _T_628 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  _T_629 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  _T_630 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  _T_631 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  _T_632 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  _T_633 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  _T_634 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  _T_635 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  _T_636 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  _T_637 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  _T_638 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  _T_639 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  _T_640 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  _T_641 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  _T_642 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  _T_643 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  _T_644 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  _T_645 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  _T_646 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  _T_647 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  _T_648 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  _T_649 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  _T_650 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  _T_651 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  _T_652 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  _T_653 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  _T_654 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  _T_655 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  _T_656 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  _T_657 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  _T_658 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  _T_659 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  _T_660 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  _T_661 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  _T_662 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  _T_663 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  _T_664 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  _T_665 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  _T_666 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  _T_667 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  _T_668 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  _T_669 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  _T_670 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  _T_671 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  _T_672 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  _T_673 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  _T_674 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  _T_675 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  _T_676 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  _T_677 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  _T_678 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  _T_679 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  _T_680 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  _T_681 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  _T_682 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  _T_683 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  _T_684 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  _T_685 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  _T_686 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  _T_687 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  _T_688 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  _T_689 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  _T_690 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  _T_691 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  _T_692 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  _T_693 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  _T_694 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  _T_695 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  _T_696 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  _T_697 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  _T_698 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  _T_699 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  _T_700 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  _T_701 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  _T_702 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  _T_703 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  _T_704 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  _T_705 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  _T_706 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  _T_707 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  _T_708 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  _T_709 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  _T_710 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  _T_711 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  _T_712 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  _T_713 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  _T_714 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  _T_715 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  _T_716 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  _T_717 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  _T_718 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  _T_719 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  _T_720 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  _T_721 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  _T_722 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  _T_723 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  _T_724 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  _T_725 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  _T_726 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  _T_727 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  _T_728 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  _T_729 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  _T_730 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  _T_731 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  _T_732 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  _T_733 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  _T_734 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  _T_735 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  _T_736 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  _T_737 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  _T_738 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  _T_739 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  _T_740 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  _T_741 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  _T_742 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  _T_743 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  _T_744 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  _T_745 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  _T_746 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  _T_747 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  _T_748 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  _T_749 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  _T_750 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  _T_751 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  _T_752 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  _T_753 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  _T_754 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  _T_755 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  _T_756 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  _T_757 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  _T_758 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  _T_759 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  _T_760 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  _T_761 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  _T_762 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  _T_763 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  _T_764 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  _T_765 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  _T_766 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  _T_767 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  _T_768 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  _T_769 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  _T_770 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  _T_771 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  _T_772 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  _T_773 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  _T_774 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  _T_775 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  _T_776 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  _T_777 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  _T_778 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  _T_779 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  _T_780 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  _T_781 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  _T_782 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  _T_783 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  _T_784 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  _T_785 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  _T_786 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  _T_787 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  _T_788 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  _T_789 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  _T_790 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  _T_791 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  _T_792 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  _T_793 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  _T_794 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  _T_795 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  _T_796 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  _T_797 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  _T_798 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  _T_799 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  _T_800 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  _T_801 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  _T_802 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  _T_803 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  _T_804 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  _T_805 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  _T_806 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  _T_807 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  _T_808 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  _T_809 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  _T_810 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  _T_811 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  _T_812 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  _T_813 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  _T_814 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  _T_815 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  _T_816 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  _T_817 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  _T_818 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  _T_819 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  _T_820 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  _T_821 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  _T_822 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  _T_823 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  _T_824 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  _T_825 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  _T_826 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  _T_827 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  _T_828 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  _T_829 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  _T_830 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  _T_831 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  _T_832 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  _T_833 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  _T_834 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  _T_835 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  _T_836 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  _T_837 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  _T_838 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  _T_839 = _RAND_773[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(rambank0_re__T_69_en & rambank0_re__T_69_mask) begin
      rambank0_re[rambank0_re__T_69_addr] <= rambank0_re__T_69_data; // @[Reorder.scala 20:21]
    end
    if(rambank0_im__T_69_en & rambank0_im__T_69_mask) begin
      rambank0_im[rambank0_im__T_69_addr] <= rambank0_im__T_69_data; // @[Reorder.scala 20:21]
    end
    if(rambank1_re__T_71_en & rambank1_re__T_71_mask) begin
      rambank1_re[rambank1_re__T_71_addr] <= rambank1_re__T_71_data; // @[Reorder.scala 21:21]
    end
    if(rambank1_im__T_71_en & rambank1_im__T_71_mask) begin
      rambank1_im[rambank1_im__T_71_addr] <= rambank1_im__T_71_data; // @[Reorder.scala 21:21]
    end
    if (reset) begin
      in_counter <= 8'h0;
    end else if (_T_65) begin
      in_counter <= _T_67;
    end
    if (reset) begin
      out_counter <= 9'h0;
    end else if (io_out_valid) begin
      out_counter <= _T_842;
    end
    _T_72 <= io_in_valid;
    _T_73 <= _T_72;
    _T_74 <= _T_73;
    _T_75 <= _T_74;
    _T_76 <= _T_75;
    _T_77 <= _T_76;
    _T_78 <= _T_77;
    _T_79 <= _T_78;
    _T_80 <= _T_79;
    _T_81 <= _T_80;
    _T_82 <= _T_81;
    _T_83 <= _T_82;
    _T_84 <= _T_83;
    _T_85 <= _T_84;
    _T_86 <= _T_85;
    _T_87 <= _T_86;
    _T_88 <= _T_87;
    _T_89 <= _T_88;
    _T_90 <= _T_89;
    _T_91 <= _T_90;
    _T_92 <= _T_91;
    _T_93 <= _T_92;
    _T_94 <= _T_93;
    _T_95 <= _T_94;
    _T_96 <= _T_95;
    _T_97 <= _T_96;
    _T_98 <= _T_97;
    _T_99 <= _T_98;
    _T_100 <= _T_99;
    _T_101 <= _T_100;
    _T_102 <= _T_101;
    _T_103 <= _T_102;
    _T_104 <= _T_103;
    _T_105 <= _T_104;
    _T_106 <= _T_105;
    _T_107 <= _T_106;
    _T_108 <= _T_107;
    _T_109 <= _T_108;
    _T_110 <= _T_109;
    _T_111 <= _T_110;
    _T_112 <= _T_111;
    _T_113 <= _T_112;
    _T_114 <= _T_113;
    _T_115 <= _T_114;
    _T_116 <= _T_115;
    _T_117 <= _T_116;
    _T_118 <= _T_117;
    _T_119 <= _T_118;
    _T_120 <= _T_119;
    _T_121 <= _T_120;
    _T_122 <= _T_121;
    _T_123 <= _T_122;
    _T_124 <= _T_123;
    _T_125 <= _T_124;
    _T_126 <= _T_125;
    _T_127 <= _T_126;
    _T_128 <= _T_127;
    _T_129 <= _T_128;
    _T_130 <= _T_129;
    _T_131 <= _T_130;
    _T_132 <= _T_131;
    _T_133 <= _T_132;
    _T_134 <= _T_133;
    _T_135 <= _T_134;
    _T_136 <= _T_135;
    _T_137 <= _T_136;
    _T_138 <= _T_137;
    _T_139 <= _T_138;
    _T_140 <= _T_139;
    _T_141 <= _T_140;
    _T_142 <= _T_141;
    _T_143 <= _T_142;
    _T_144 <= _T_143;
    _T_145 <= _T_144;
    _T_146 <= _T_145;
    _T_147 <= _T_146;
    _T_148 <= _T_147;
    _T_149 <= _T_148;
    _T_150 <= _T_149;
    _T_151 <= _T_150;
    _T_152 <= _T_151;
    _T_153 <= _T_152;
    _T_154 <= _T_153;
    _T_155 <= _T_154;
    _T_156 <= _T_155;
    _T_157 <= _T_156;
    _T_158 <= _T_157;
    _T_159 <= _T_158;
    _T_160 <= _T_159;
    _T_161 <= _T_160;
    _T_162 <= _T_161;
    _T_163 <= _T_162;
    _T_164 <= _T_163;
    _T_165 <= _T_164;
    _T_166 <= _T_165;
    _T_167 <= _T_166;
    _T_168 <= _T_167;
    _T_169 <= _T_168;
    _T_170 <= _T_169;
    _T_171 <= _T_170;
    _T_172 <= _T_171;
    _T_173 <= _T_172;
    _T_174 <= _T_173;
    _T_175 <= _T_174;
    _T_176 <= _T_175;
    _T_177 <= _T_176;
    _T_178 <= _T_177;
    _T_179 <= _T_178;
    _T_180 <= _T_179;
    _T_181 <= _T_180;
    _T_182 <= _T_181;
    _T_183 <= _T_182;
    _T_184 <= _T_183;
    _T_185 <= _T_184;
    _T_186 <= _T_185;
    _T_187 <= _T_186;
    _T_188 <= _T_187;
    _T_189 <= _T_188;
    _T_190 <= _T_189;
    _T_191 <= _T_190;
    _T_192 <= _T_191;
    _T_193 <= _T_192;
    _T_194 <= _T_193;
    _T_195 <= _T_194;
    _T_196 <= _T_195;
    _T_197 <= _T_196;
    _T_198 <= _T_197;
    _T_199 <= _T_198;
    _T_200 <= _T_199;
    _T_201 <= _T_200;
    _T_202 <= _T_201;
    _T_203 <= _T_202;
    _T_204 <= _T_203;
    _T_205 <= _T_204;
    _T_206 <= _T_205;
    _T_207 <= _T_206;
    _T_208 <= _T_207;
    _T_209 <= _T_208;
    _T_210 <= _T_209;
    _T_211 <= _T_210;
    _T_212 <= _T_211;
    _T_213 <= _T_212;
    _T_214 <= _T_213;
    _T_215 <= _T_214;
    _T_216 <= _T_215;
    _T_217 <= _T_216;
    _T_218 <= _T_217;
    _T_219 <= _T_218;
    _T_220 <= _T_219;
    _T_221 <= _T_220;
    _T_222 <= _T_221;
    _T_223 <= _T_222;
    _T_224 <= _T_223;
    _T_225 <= _T_224;
    _T_226 <= _T_225;
    _T_227 <= _T_226;
    _T_228 <= _T_227;
    _T_229 <= _T_228;
    _T_230 <= _T_229;
    _T_231 <= _T_230;
    _T_232 <= _T_231;
    _T_233 <= _T_232;
    _T_234 <= _T_233;
    _T_235 <= _T_234;
    _T_236 <= _T_235;
    _T_237 <= _T_236;
    _T_238 <= _T_237;
    _T_239 <= _T_238;
    _T_240 <= _T_239;
    _T_241 <= _T_240;
    _T_242 <= _T_241;
    _T_243 <= _T_242;
    _T_244 <= _T_243;
    _T_245 <= _T_244;
    _T_246 <= _T_245;
    _T_247 <= _T_246;
    _T_248 <= _T_247;
    _T_249 <= _T_248;
    _T_250 <= _T_249;
    _T_251 <= _T_250;
    _T_252 <= _T_251;
    _T_253 <= _T_252;
    _T_254 <= _T_253;
    _T_255 <= _T_254;
    _T_256 <= _T_255;
    _T_257 <= _T_256;
    _T_258 <= _T_257;
    _T_259 <= _T_258;
    _T_260 <= _T_259;
    _T_261 <= _T_260;
    _T_262 <= _T_261;
    _T_263 <= _T_262;
    _T_264 <= _T_263;
    _T_265 <= _T_264;
    _T_266 <= _T_265;
    _T_267 <= _T_266;
    _T_268 <= _T_267;
    _T_269 <= _T_268;
    _T_270 <= _T_269;
    _T_271 <= _T_270;
    _T_272 <= _T_271;
    _T_273 <= _T_272;
    _T_274 <= _T_273;
    _T_275 <= _T_274;
    _T_276 <= _T_275;
    _T_277 <= _T_276;
    _T_278 <= _T_277;
    _T_279 <= _T_278;
    _T_280 <= _T_279;
    _T_281 <= _T_280;
    _T_282 <= _T_281;
    _T_283 <= _T_282;
    _T_284 <= _T_283;
    _T_285 <= _T_284;
    _T_286 <= _T_285;
    _T_287 <= _T_286;
    _T_288 <= _T_287;
    _T_289 <= _T_288;
    _T_290 <= _T_289;
    _T_291 <= _T_290;
    _T_292 <= _T_291;
    _T_293 <= _T_292;
    _T_294 <= _T_293;
    _T_295 <= _T_294;
    _T_296 <= _T_295;
    _T_297 <= _T_296;
    _T_298 <= _T_297;
    _T_299 <= _T_298;
    _T_300 <= _T_299;
    _T_301 <= _T_300;
    _T_302 <= _T_301;
    _T_303 <= _T_302;
    _T_304 <= _T_303;
    _T_305 <= _T_304;
    _T_306 <= _T_305;
    _T_307 <= _T_306;
    _T_308 <= _T_307;
    _T_309 <= _T_308;
    _T_310 <= _T_309;
    _T_311 <= _T_310;
    _T_312 <= _T_311;
    _T_313 <= _T_312;
    _T_314 <= _T_313;
    _T_315 <= _T_314;
    _T_316 <= _T_315;
    _T_317 <= _T_316;
    _T_318 <= _T_317;
    _T_319 <= _T_318;
    _T_320 <= _T_319;
    _T_321 <= _T_320;
    _T_322 <= _T_321;
    _T_323 <= _T_322;
    _T_324 <= _T_323;
    _T_325 <= _T_324;
    _T_326 <= _T_325;
    _T_327 <= _T_326;
    _T_328 <= io_in_valid;
    _T_329 <= _T_328;
    _T_330 <= _T_329;
    _T_331 <= _T_330;
    _T_332 <= _T_331;
    _T_333 <= _T_332;
    _T_334 <= _T_333;
    _T_335 <= _T_334;
    _T_336 <= _T_335;
    _T_337 <= _T_336;
    _T_338 <= _T_337;
    _T_339 <= _T_338;
    _T_340 <= _T_339;
    _T_341 <= _T_340;
    _T_342 <= _T_341;
    _T_343 <= _T_342;
    _T_344 <= _T_343;
    _T_345 <= _T_344;
    _T_346 <= _T_345;
    _T_347 <= _T_346;
    _T_348 <= _T_347;
    _T_349 <= _T_348;
    _T_350 <= _T_349;
    _T_351 <= _T_350;
    _T_352 <= _T_351;
    _T_353 <= _T_352;
    _T_354 <= _T_353;
    _T_355 <= _T_354;
    _T_356 <= _T_355;
    _T_357 <= _T_356;
    _T_358 <= _T_357;
    _T_359 <= _T_358;
    _T_360 <= _T_359;
    _T_361 <= _T_360;
    _T_362 <= _T_361;
    _T_363 <= _T_362;
    _T_364 <= _T_363;
    _T_365 <= _T_364;
    _T_366 <= _T_365;
    _T_367 <= _T_366;
    _T_368 <= _T_367;
    _T_369 <= _T_368;
    _T_370 <= _T_369;
    _T_371 <= _T_370;
    _T_372 <= _T_371;
    _T_373 <= _T_372;
    _T_374 <= _T_373;
    _T_375 <= _T_374;
    _T_376 <= _T_375;
    _T_377 <= _T_376;
    _T_378 <= _T_377;
    _T_379 <= _T_378;
    _T_380 <= _T_379;
    _T_381 <= _T_380;
    _T_382 <= _T_381;
    _T_383 <= _T_382;
    _T_384 <= _T_383;
    _T_385 <= _T_384;
    _T_386 <= _T_385;
    _T_387 <= _T_386;
    _T_388 <= _T_387;
    _T_389 <= _T_388;
    _T_390 <= _T_389;
    _T_391 <= _T_390;
    _T_392 <= _T_391;
    _T_393 <= _T_392;
    _T_394 <= _T_393;
    _T_395 <= _T_394;
    _T_396 <= _T_395;
    _T_397 <= _T_396;
    _T_398 <= _T_397;
    _T_399 <= _T_398;
    _T_400 <= _T_399;
    _T_401 <= _T_400;
    _T_402 <= _T_401;
    _T_403 <= _T_402;
    _T_404 <= _T_403;
    _T_405 <= _T_404;
    _T_406 <= _T_405;
    _T_407 <= _T_406;
    _T_408 <= _T_407;
    _T_409 <= _T_408;
    _T_410 <= _T_409;
    _T_411 <= _T_410;
    _T_412 <= _T_411;
    _T_413 <= _T_412;
    _T_414 <= _T_413;
    _T_415 <= _T_414;
    _T_416 <= _T_415;
    _T_417 <= _T_416;
    _T_418 <= _T_417;
    _T_419 <= _T_418;
    _T_420 <= _T_419;
    _T_421 <= _T_420;
    _T_422 <= _T_421;
    _T_423 <= _T_422;
    _T_424 <= _T_423;
    _T_425 <= _T_424;
    _T_426 <= _T_425;
    _T_427 <= _T_426;
    _T_428 <= _T_427;
    _T_429 <= _T_428;
    _T_430 <= _T_429;
    _T_431 <= _T_430;
    _T_432 <= _T_431;
    _T_433 <= _T_432;
    _T_434 <= _T_433;
    _T_435 <= _T_434;
    _T_436 <= _T_435;
    _T_437 <= _T_436;
    _T_438 <= _T_437;
    _T_439 <= _T_438;
    _T_440 <= _T_439;
    _T_441 <= _T_440;
    _T_442 <= _T_441;
    _T_443 <= _T_442;
    _T_444 <= _T_443;
    _T_445 <= _T_444;
    _T_446 <= _T_445;
    _T_447 <= _T_446;
    _T_448 <= _T_447;
    _T_449 <= _T_448;
    _T_450 <= _T_449;
    _T_451 <= _T_450;
    _T_452 <= _T_451;
    _T_453 <= _T_452;
    _T_454 <= _T_453;
    _T_455 <= _T_454;
    _T_456 <= _T_455;
    _T_457 <= _T_456;
    _T_458 <= _T_457;
    _T_459 <= _T_458;
    _T_460 <= _T_459;
    _T_461 <= _T_460;
    _T_462 <= _T_461;
    _T_463 <= _T_462;
    _T_464 <= _T_463;
    _T_465 <= _T_464;
    _T_466 <= _T_465;
    _T_467 <= _T_466;
    _T_468 <= _T_467;
    _T_469 <= _T_468;
    _T_470 <= _T_469;
    _T_471 <= _T_470;
    _T_472 <= _T_471;
    _T_473 <= _T_472;
    _T_474 <= _T_473;
    _T_475 <= _T_474;
    _T_476 <= _T_475;
    _T_477 <= _T_476;
    _T_478 <= _T_477;
    _T_479 <= _T_478;
    _T_480 <= _T_479;
    _T_481 <= _T_480;
    _T_482 <= _T_481;
    _T_483 <= _T_482;
    _T_484 <= _T_483;
    _T_485 <= _T_484;
    _T_486 <= _T_485;
    _T_487 <= _T_486;
    _T_488 <= _T_487;
    _T_489 <= _T_488;
    _T_490 <= _T_489;
    _T_491 <= _T_490;
    _T_492 <= _T_491;
    _T_493 <= _T_492;
    _T_494 <= _T_493;
    _T_495 <= _T_494;
    _T_496 <= _T_495;
    _T_497 <= _T_496;
    _T_498 <= _T_497;
    _T_499 <= _T_498;
    _T_500 <= _T_499;
    _T_501 <= _T_500;
    _T_502 <= _T_501;
    _T_503 <= _T_502;
    _T_504 <= _T_503;
    _T_505 <= _T_504;
    _T_506 <= _T_505;
    _T_507 <= _T_506;
    _T_508 <= _T_507;
    _T_509 <= _T_508;
    _T_510 <= _T_509;
    _T_511 <= _T_510;
    _T_512 <= _T_511;
    _T_513 <= _T_512;
    _T_514 <= _T_513;
    _T_515 <= _T_514;
    _T_516 <= _T_515;
    _T_517 <= _T_516;
    _T_518 <= _T_517;
    _T_519 <= _T_518;
    _T_520 <= _T_519;
    _T_521 <= _T_520;
    _T_522 <= _T_521;
    _T_523 <= _T_522;
    _T_524 <= _T_523;
    _T_525 <= _T_524;
    _T_526 <= _T_525;
    _T_527 <= _T_526;
    _T_528 <= _T_527;
    _T_529 <= _T_528;
    _T_530 <= _T_529;
    _T_531 <= _T_530;
    _T_532 <= _T_531;
    _T_533 <= _T_532;
    _T_534 <= _T_533;
    _T_535 <= _T_534;
    _T_536 <= _T_535;
    _T_537 <= _T_536;
    _T_538 <= _T_537;
    _T_539 <= _T_538;
    _T_540 <= _T_539;
    _T_541 <= _T_540;
    _T_542 <= _T_541;
    _T_543 <= _T_542;
    _T_544 <= _T_543;
    _T_545 <= _T_544;
    _T_546 <= _T_545;
    _T_547 <= _T_546;
    _T_548 <= _T_547;
    _T_549 <= _T_548;
    _T_550 <= _T_549;
    _T_551 <= _T_550;
    _T_552 <= _T_551;
    _T_553 <= _T_552;
    _T_554 <= _T_553;
    _T_555 <= _T_554;
    _T_556 <= _T_555;
    _T_557 <= _T_556;
    _T_558 <= _T_557;
    _T_559 <= _T_558;
    _T_560 <= _T_559;
    _T_561 <= _T_560;
    _T_562 <= _T_561;
    _T_563 <= _T_562;
    _T_564 <= _T_563;
    _T_565 <= _T_564;
    _T_566 <= _T_565;
    _T_567 <= _T_566;
    _T_568 <= _T_567;
    _T_569 <= _T_568;
    _T_570 <= _T_569;
    _T_571 <= _T_570;
    _T_572 <= _T_571;
    _T_573 <= _T_572;
    _T_574 <= _T_573;
    _T_575 <= _T_574;
    _T_576 <= _T_575;
    _T_577 <= _T_576;
    _T_578 <= _T_577;
    _T_579 <= _T_578;
    _T_580 <= _T_579;
    _T_581 <= _T_580;
    _T_582 <= _T_581;
    _T_583 <= _T_582;
    _T_584 <= _T_583;
    _T_585 <= _T_584;
    _T_586 <= _T_585;
    _T_587 <= _T_586;
    _T_588 <= _T_587;
    _T_589 <= _T_588;
    _T_590 <= _T_589;
    _T_591 <= _T_590;
    _T_592 <= _T_591;
    _T_593 <= _T_592;
    _T_594 <= _T_593;
    _T_595 <= _T_594;
    _T_596 <= _T_595;
    _T_597 <= _T_596;
    _T_598 <= _T_597;
    _T_599 <= _T_598;
    _T_600 <= _T_599;
    _T_601 <= _T_600;
    _T_602 <= _T_601;
    _T_603 <= _T_602;
    _T_604 <= _T_603;
    _T_605 <= _T_604;
    _T_606 <= _T_605;
    _T_607 <= _T_606;
    _T_608 <= _T_607;
    _T_609 <= _T_608;
    _T_610 <= _T_609;
    _T_611 <= _T_610;
    _T_612 <= _T_611;
    _T_613 <= _T_612;
    _T_614 <= _T_613;
    _T_615 <= _T_614;
    _T_616 <= _T_615;
    _T_617 <= _T_616;
    _T_618 <= _T_617;
    _T_619 <= _T_618;
    _T_620 <= _T_619;
    _T_621 <= _T_620;
    _T_622 <= _T_621;
    _T_623 <= _T_622;
    _T_624 <= _T_623;
    _T_625 <= _T_624;
    _T_626 <= _T_625;
    _T_627 <= _T_626;
    _T_628 <= _T_627;
    _T_629 <= _T_628;
    _T_630 <= _T_629;
    _T_631 <= _T_630;
    _T_632 <= _T_631;
    _T_633 <= _T_632;
    _T_634 <= _T_633;
    _T_635 <= _T_634;
    _T_636 <= _T_635;
    _T_637 <= _T_636;
    _T_638 <= _T_637;
    _T_639 <= _T_638;
    _T_640 <= _T_639;
    _T_641 <= _T_640;
    _T_642 <= _T_641;
    _T_643 <= _T_642;
    _T_644 <= _T_643;
    _T_645 <= _T_644;
    _T_646 <= _T_645;
    _T_647 <= _T_646;
    _T_648 <= _T_647;
    _T_649 <= _T_648;
    _T_650 <= _T_649;
    _T_651 <= _T_650;
    _T_652 <= _T_651;
    _T_653 <= _T_652;
    _T_654 <= _T_653;
    _T_655 <= _T_654;
    _T_656 <= _T_655;
    _T_657 <= _T_656;
    _T_658 <= _T_657;
    _T_659 <= _T_658;
    _T_660 <= _T_659;
    _T_661 <= _T_660;
    _T_662 <= _T_661;
    _T_663 <= _T_662;
    _T_664 <= _T_663;
    _T_665 <= _T_664;
    _T_666 <= _T_665;
    _T_667 <= _T_666;
    _T_668 <= _T_667;
    _T_669 <= _T_668;
    _T_670 <= _T_669;
    _T_671 <= _T_670;
    _T_672 <= _T_671;
    _T_673 <= _T_672;
    _T_674 <= _T_673;
    _T_675 <= _T_674;
    _T_676 <= _T_675;
    _T_677 <= _T_676;
    _T_678 <= _T_677;
    _T_679 <= _T_678;
    _T_680 <= _T_679;
    _T_681 <= _T_680;
    _T_682 <= _T_681;
    _T_683 <= _T_682;
    _T_684 <= _T_683;
    _T_685 <= _T_684;
    _T_686 <= _T_685;
    _T_687 <= _T_686;
    _T_688 <= _T_687;
    _T_689 <= _T_688;
    _T_690 <= _T_689;
    _T_691 <= _T_690;
    _T_692 <= _T_691;
    _T_693 <= _T_692;
    _T_694 <= _T_693;
    _T_695 <= _T_694;
    _T_696 <= _T_695;
    _T_697 <= _T_696;
    _T_698 <= _T_697;
    _T_699 <= _T_698;
    _T_700 <= _T_699;
    _T_701 <= _T_700;
    _T_702 <= _T_701;
    _T_703 <= _T_702;
    _T_704 <= _T_703;
    _T_705 <= _T_704;
    _T_706 <= _T_705;
    _T_707 <= _T_706;
    _T_708 <= _T_707;
    _T_709 <= _T_708;
    _T_710 <= _T_709;
    _T_711 <= _T_710;
    _T_712 <= _T_711;
    _T_713 <= _T_712;
    _T_714 <= _T_713;
    _T_715 <= _T_714;
    _T_716 <= _T_715;
    _T_717 <= _T_716;
    _T_718 <= _T_717;
    _T_719 <= _T_718;
    _T_720 <= _T_719;
    _T_721 <= _T_720;
    _T_722 <= _T_721;
    _T_723 <= _T_722;
    _T_724 <= _T_723;
    _T_725 <= _T_724;
    _T_726 <= _T_725;
    _T_727 <= _T_726;
    _T_728 <= _T_727;
    _T_729 <= _T_728;
    _T_730 <= _T_729;
    _T_731 <= _T_730;
    _T_732 <= _T_731;
    _T_733 <= _T_732;
    _T_734 <= _T_733;
    _T_735 <= _T_734;
    _T_736 <= _T_735;
    _T_737 <= _T_736;
    _T_738 <= _T_737;
    _T_739 <= _T_738;
    _T_740 <= _T_739;
    _T_741 <= _T_740;
    _T_742 <= _T_741;
    _T_743 <= _T_742;
    _T_744 <= _T_743;
    _T_745 <= _T_744;
    _T_746 <= _T_745;
    _T_747 <= _T_746;
    _T_748 <= _T_747;
    _T_749 <= _T_748;
    _T_750 <= _T_749;
    _T_751 <= _T_750;
    _T_752 <= _T_751;
    _T_753 <= _T_752;
    _T_754 <= _T_753;
    _T_755 <= _T_754;
    _T_756 <= _T_755;
    _T_757 <= _T_756;
    _T_758 <= _T_757;
    _T_759 <= _T_758;
    _T_760 <= _T_759;
    _T_761 <= _T_760;
    _T_762 <= _T_761;
    _T_763 <= _T_762;
    _T_764 <= _T_763;
    _T_765 <= _T_764;
    _T_766 <= _T_765;
    _T_767 <= _T_766;
    _T_768 <= _T_767;
    _T_769 <= _T_768;
    _T_770 <= _T_769;
    _T_771 <= _T_770;
    _T_772 <= _T_771;
    _T_773 <= _T_772;
    _T_774 <= _T_773;
    _T_775 <= _T_774;
    _T_776 <= _T_775;
    _T_777 <= _T_776;
    _T_778 <= _T_777;
    _T_779 <= _T_778;
    _T_780 <= _T_779;
    _T_781 <= _T_780;
    _T_782 <= _T_781;
    _T_783 <= _T_782;
    _T_784 <= _T_783;
    _T_785 <= _T_784;
    _T_786 <= _T_785;
    _T_787 <= _T_786;
    _T_788 <= _T_787;
    _T_789 <= _T_788;
    _T_790 <= _T_789;
    _T_791 <= _T_790;
    _T_792 <= _T_791;
    _T_793 <= _T_792;
    _T_794 <= _T_793;
    _T_795 <= _T_794;
    _T_796 <= _T_795;
    _T_797 <= _T_796;
    _T_798 <= _T_797;
    _T_799 <= _T_798;
    _T_800 <= _T_799;
    _T_801 <= _T_800;
    _T_802 <= _T_801;
    _T_803 <= _T_802;
    _T_804 <= _T_803;
    _T_805 <= _T_804;
    _T_806 <= _T_805;
    _T_807 <= _T_806;
    _T_808 <= _T_807;
    _T_809 <= _T_808;
    _T_810 <= _T_809;
    _T_811 <= _T_810;
    _T_812 <= _T_811;
    _T_813 <= _T_812;
    _T_814 <= _T_813;
    _T_815 <= _T_814;
    _T_816 <= _T_815;
    _T_817 <= _T_816;
    _T_818 <= _T_817;
    _T_819 <= _T_818;
    _T_820 <= _T_819;
    _T_821 <= _T_820;
    _T_822 <= _T_821;
    _T_823 <= _T_822;
    _T_824 <= _T_823;
    _T_825 <= _T_824;
    _T_826 <= _T_825;
    _T_827 <= _T_826;
    _T_828 <= _T_827;
    _T_829 <= _T_828;
    _T_830 <= _T_829;
    _T_831 <= _T_830;
    _T_832 <= _T_831;
    _T_833 <= _T_832;
    _T_834 <= _T_833;
    _T_835 <= _T_834;
    _T_836 <= _T_835;
    _T_837 <= _T_836;
    _T_838 <= _T_837;
    _T_839 <= _T_838;
  end
endmodule
module FFTReorder(
  input         clock,
  input         reset,
  input  [31:0] io_dIn_re,
  input  [31:0] io_dIn_im,
  input         io_din_valid,
  output [31:0] io_dOut_re,
  output [31:0] io_dOut_im,
  output        io_dout_valid
);
  wire  fftblock_clock; // @[Reorder.scala 62:29]
  wire  fftblock_reset; // @[Reorder.scala 62:29]
  wire [31:0] fftblock_io_dIn_re; // @[Reorder.scala 62:29]
  wire [31:0] fftblock_io_dIn_im; // @[Reorder.scala 62:29]
  wire  fftblock_io_din_valid; // @[Reorder.scala 62:29]
  wire [31:0] fftblock_io_dOut1_re; // @[Reorder.scala 62:29]
  wire [31:0] fftblock_io_dOut1_im; // @[Reorder.scala 62:29]
  wire [31:0] fftblock_io_dOut2_re; // @[Reorder.scala 62:29]
  wire [31:0] fftblock_io_dOut2_im; // @[Reorder.scala 62:29]
  wire  fftblock_io_dout_valid; // @[Reorder.scala 62:29]
  wire  reorderblock_clock; // @[Reorder.scala 66:28]
  wire  reorderblock_reset; // @[Reorder.scala 66:28]
  wire [31:0] reorderblock_io_in1_re; // @[Reorder.scala 66:28]
  wire [31:0] reorderblock_io_in1_im; // @[Reorder.scala 66:28]
  wire [31:0] reorderblock_io_in2_re; // @[Reorder.scala 66:28]
  wire [31:0] reorderblock_io_in2_im; // @[Reorder.scala 66:28]
  wire  reorderblock_io_in_valid; // @[Reorder.scala 66:28]
  wire [31:0] reorderblock_io_out_re; // @[Reorder.scala 66:28]
  wire [31:0] reorderblock_io_out_im; // @[Reorder.scala 66:28]
  wire  reorderblock_io_out_valid; // @[Reorder.scala 66:28]
  FFT fftblock ( // @[Reorder.scala 62:29]
    .clock(fftblock_clock),
    .reset(fftblock_reset),
    .io_dIn_re(fftblock_io_dIn_re),
    .io_dIn_im(fftblock_io_dIn_im),
    .io_din_valid(fftblock_io_din_valid),
    .io_dOut1_re(fftblock_io_dOut1_re),
    .io_dOut1_im(fftblock_io_dOut1_im),
    .io_dOut2_re(fftblock_io_dOut2_re),
    .io_dOut2_im(fftblock_io_dOut2_im),
    .io_dout_valid(fftblock_io_dout_valid)
  );
  Reorder reorderblock ( // @[Reorder.scala 66:28]
    .clock(reorderblock_clock),
    .reset(reorderblock_reset),
    .io_in1_re(reorderblock_io_in1_re),
    .io_in1_im(reorderblock_io_in1_im),
    .io_in2_re(reorderblock_io_in2_re),
    .io_in2_im(reorderblock_io_in2_im),
    .io_in_valid(reorderblock_io_in_valid),
    .io_out_re(reorderblock_io_out_re),
    .io_out_im(reorderblock_io_out_im),
    .io_out_valid(reorderblock_io_out_valid)
  );
  assign io_dOut_re = reorderblock_io_out_re; // @[Reorder.scala 71:11]
  assign io_dOut_im = reorderblock_io_out_im; // @[Reorder.scala 71:11]
  assign io_dout_valid = reorderblock_io_out_valid; // @[Reorder.scala 72:17]
  assign fftblock_clock = clock;
  assign fftblock_reset = reset;
  assign fftblock_io_dIn_re = io_dIn_re; // @[Reorder.scala 63:19]
  assign fftblock_io_dIn_im = io_dIn_im; // @[Reorder.scala 63:19]
  assign fftblock_io_din_valid = io_din_valid; // @[Reorder.scala 64:25]
  assign reorderblock_clock = clock;
  assign reorderblock_reset = reset;
  assign reorderblock_io_in1_re = fftblock_io_dOut1_re; // @[Reorder.scala 67:23]
  assign reorderblock_io_in1_im = fftblock_io_dOut1_im; // @[Reorder.scala 67:23]
  assign reorderblock_io_in2_re = fftblock_io_dOut2_re; // @[Reorder.scala 68:23]
  assign reorderblock_io_in2_im = fftblock_io_dOut2_im; // @[Reorder.scala 68:23]
  assign reorderblock_io_in_valid = fftblock_io_dout_valid; // @[Reorder.scala 69:28]
endmodule
